* NGSPICE file created from uart_macro_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

.subckt uart_macro_wrapper io_oeb[0] io_oeb[1] uart_irq uart_rx uart_tx vccd1 vssd1
+ wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3155_ _3579_/CLK _3155_/D vssd1 vssd1 vccd1 vccd1 _3155_/Q sky130_fd_sc_hd__dfxtp_1
X_2106_ _2079_/X _2106_/B vssd1 vssd1 vccd1 vccd1 _2106_/X sky130_fd_sc_hd__and2b_1
X_3086_ _3090_/A vssd1 vssd1 vccd1 vccd1 _3086_/Y sky130_fd_sc_hd__inv_2
X_2037_ hold142/X _3281_/Q _3272_/Q _3263_/Q _2221_/B _2219_/A vssd1 vssd1 vccd1 vccd1
+ _2037_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2651__A0 _2360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2939_ _3127_/A vssd1 vssd1 vccd1 vccd1 _2939_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_72_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold340 _2753_/X vssd1 vssd1 vccd1 vccd1 _3282_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold362 _1620_/X vssd1 vssd1 vccd1 vccd1 _3636_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 _3293_/Q vssd1 vssd1 vccd1 vccd1 hold351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 _2793_/X vssd1 vssd1 vccd1 vccd1 _3318_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 _3304_/Q vssd1 vssd1 vccd1 vccd1 hold384/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold395 _2694_/X vssd1 vssd1 vccd1 vccd1 _3231_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 _3568_/Q vssd1 vssd1 vccd1 vccd1 hold786/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1040 _3625_/Q vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2642__A0 _2355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1684__A1 _2401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2633__A0 _2356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__1610__C input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2724_ _2805_/A1 hold386/X _2728_/S vssd1 vssd1 vccd1 vccd1 _2724_/X sky130_fd_sc_hd__mux2_1
X_2655_ _3487_/Q hold36/X _3488_/Q vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__nand3b_1
X_1606_ _1607_/A _1607_/B vssd1 vssd1 vccd1 vccd1 _2577_/B sky130_fd_sc_hd__and2_1
XFILLER_0_1_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2586_ hold447/X _2806_/A1 _2589_/S vssd1 vssd1 vccd1 vccd1 _2586_/X sky130_fd_sc_hd__mux2_1
Xfanout127 _3057_/A vssd1 vssd1 vccd1 vccd1 _3032_/A sky130_fd_sc_hd__buf_8
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout116 _3112_/A vssd1 vssd1 vccd1 vccd1 _3069_/A sky130_fd_sc_hd__buf_6
Xfanout105 hold75/X vssd1 vssd1 vccd1 vccd1 _2805_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2884__S _2890_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3207_ _3333_/CLK _3207_/D vssd1 vssd1 vccd1 vccd1 _3207_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2872__A0 _2358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3138_ _3333_/CLK _3138_/D vssd1 vssd1 vccd1 vccd1 _3138_/Q sky130_fd_sc_hd__dfxtp_1
X_3069_ _3069_/A vssd1 vssd1 vccd1 vccd1 _3069_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold170 _2794_/X vssd1 vssd1 vccd1 vccd1 _3319_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _3612_/Q vssd1 vssd1 vccd1 vccd1 _1570_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 _3242_/Q vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2794__S _2799_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2615__A0 _2358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3654__A _3655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2440_ _3480_/Q _2507_/B _2508_/A vssd1 vssd1 vccd1 vccd1 _2440_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2371_ hold940/X _2377_/C _2370_/Y _2144_/D vssd1 vssd1 vccd1 vccd1 _2371_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2529__S0 _2532_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2854__A0 _2109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2606__A0 _2109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout125_A _3057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2879__S _2880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2707_ _2406_/A hold437/X _2707_/S vssd1 vssd1 vccd1 vccd1 _2707_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2638_ _2105_/A hold726/X _2643_/S vssd1 vssd1 vccd1 vccd1 _2638_/X sky130_fd_sc_hd__mux2_1
X_2569_ _3453_/Q _2510_/B _2559_/X _2568_/X vssd1 vssd1 vccd1 vccd1 _2570_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1991__S1 _2045_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2845__A0 _2104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1648__A1 hold87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2789__S hold38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2836__A0 _2360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1639__A1 _2401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3649__A _3655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1940_ _1927_/Y _1935_/Y _1939_/X _1935_/B _2349_/B vssd1 vssd1 vccd1 vccd1 _1940_/X
+ sky130_fd_sc_hd__a32o_1
X_1871_ _1871_/A _1871_/B vssd1 vssd1 vccd1 vccd1 _1871_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1811__A1 _2383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3610_ _3610_/CLK _3610_/D _3101_/Y vssd1 vssd1 vccd1 vccd1 _3610_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3541_ _3573_/CLK _3541_/D _3035_/Y vssd1 vssd1 vccd1 vccd1 _3541_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2699__S _2707_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold906 _3457_/Q vssd1 vssd1 vccd1 vccd1 _2270_/A sky130_fd_sc_hd__buf_1
Xhold928 _1878_/X vssd1 vssd1 vccd1 vccd1 _3527_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 _1876_/X vssd1 vssd1 vccd1 vccd1 _3528_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold939 _2156_/X vssd1 vssd1 vccd1 vccd1 _3493_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3472_ _3590_/CLK _3472_/D _2966_/Y vssd1 vssd1 vccd1 vccd1 _3472_/Q sky130_fd_sc_hd__dfstp_1
X_2423_ _3611_/Q hold52/A _2507_/C _3511_/Q vssd1 vssd1 vccd1 vccd1 _2423_/X sky130_fd_sc_hd__o22a_1
X_2354_ _2352_/X _2353_/X hold882/X vssd1 vssd1 vccd1 vccd1 _2354_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__1973__S1 _2195_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2285_ hold92/X hold50/X hold8/X _1623_/C vssd1 vssd1 vccd1 vccd1 _2413_/B sky130_fd_sc_hd__or4b_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2357__B _2357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2294__A1 hold78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2070_ _2070_/A _2096_/B vssd1 vssd1 vccd1 vccd1 _2070_/X sky130_fd_sc_hd__and2_1
XFILLER_0_72_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2972_ _3097_/A vssd1 vssd1 vccd1 vccd1 _2972_/Y sky130_fd_sc_hd__inv_2
X_1923_ _1923_/A _2162_/B _2363_/A vssd1 vssd1 vccd1 vccd1 _1932_/B sky130_fd_sc_hd__or3b_4
XFILLER_0_44_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1854_ _1837_/Y _1853_/X _1557_/A vssd1 vssd1 vccd1 vccd1 _1858_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold703 _2637_/X vssd1 vssd1 vccd1 vccd1 _3183_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1785_ _2070_/A _2092_/A _3622_/Q vssd1 vssd1 vccd1 vccd1 _1785_/Y sky130_fd_sc_hd__o21ai_2
X_3524_ _3576_/CLK _3524_/D _3018_/Y vssd1 vssd1 vccd1 vccd1 _3524_/Q sky130_fd_sc_hd__dfrtp_1
Xhold725 _2902_/X vssd1 vssd1 vccd1 vccd1 _3430_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 _3156_/Q vssd1 vssd1 vccd1 vccd1 hold714/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 _3416_/Q vssd1 vssd1 vccd1 vccd1 hold736/X sky130_fd_sc_hd__dlygate4sd3_1
X_3455_ _3633_/CLK hold57/X _2949_/Y vssd1 vssd1 vccd1 vccd1 _3455_/Q sky130_fd_sc_hd__dfrtp_1
Xhold769 _2831_/X vssd1 vssd1 vccd1 vccd1 _3362_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 _2636_/X vssd1 vssd1 vccd1 vccd1 _3182_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 _3403_/Q vssd1 vssd1 vccd1 vccd1 hold758/X sky130_fd_sc_hd__dlygate4sd3_1
X_2406_ _2406_/A hold98/X hold95/X vssd1 vssd1 vccd1 vccd1 _3588_/D sky130_fd_sc_hd__and3_1
X_3386_ _3431_/CLK _3386_/D vssd1 vssd1 vccd1 vccd1 _3386_/Q sky130_fd_sc_hd__dfxtp_1
X_2337_ _3576_/Q _2363_/A _3380_/Q vssd1 vssd1 vccd1 vccd1 _2338_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2268_ _2363_/A _2267_/X _2270_/C vssd1 vssd1 vccd1 vccd1 _2283_/A sky130_fd_sc_hd__o21a_1
XANTENNA__2892__S _2900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2199_ _2211_/A _2183_/Y _2208_/B _2184_/X vssd1 vssd1 vccd1 vccd1 _2211_/B sky130_fd_sc_hd__o31ai_4
XFILLER_0_79_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2132__S _2144_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1971__S _2036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__clkbuf_4
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2019__A1 _2036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3484_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2550__B hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1570_ _1570_/A vssd1 vssd1 vccd1 vccd1 _1570_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_34_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _3326_/CLK _3240_/D vssd1 vssd1 vccd1 vccd1 _3240_/Q sky130_fd_sc_hd__dfxtp_1
X_3171_ _3432_/CLK _3171_/D vssd1 vssd1 vccd1 vccd1 _3171_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2122_ _3497_/Q _2122_/B vssd1 vssd1 vccd1 vccd1 _2123_/D sky130_fd_sc_hd__xor2_1
XFILLER_0_83_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2053_ _2053_/A _2144_/C vssd1 vssd1 vccd1 vccd1 _2053_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2955_ _3122_/A vssd1 vssd1 vccd1 vccd1 _2955_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2886_ _2104_/B hold736/X _2890_/S vssd1 vssd1 vccd1 vccd1 _2886_/X sky130_fd_sc_hd__mux2_1
X_1906_ hold35/X _2421_/B vssd1 vssd1 vccd1 vccd1 _1908_/D sky130_fd_sc_hd__and2_2
X_1837_ _1837_/A vssd1 vssd1 vccd1 vccd1 _1837_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold511 _2822_/X vssd1 vssd1 vccd1 vccd1 _3354_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold500 _3359_/Q vssd1 vssd1 vccd1 vccd1 hold500/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 _3369_/Q vssd1 vssd1 vccd1 vccd1 hold522/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2887__S _2890_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold544 _3339_/Q vssd1 vssd1 vccd1 vccd1 hold544/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 _2609_/X vssd1 vssd1 vccd1 vccd1 _3159_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3507_ _3509_/CLK _3507_/D _3001_/Y vssd1 vssd1 vccd1 vccd1 _3507_/Q sky130_fd_sc_hd__dfrtp_1
X_1768_ _1767_/X hold929/X _1768_/S vssd1 vssd1 vccd1 vccd1 _2383_/B sky130_fd_sc_hd__mux2_4
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold588 _3336_/Q vssd1 vssd1 vccd1 vccd1 hold588/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 _2621_/X vssd1 vssd1 vccd1 vccd1 _3169_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 _3419_/Q vssd1 vssd1 vccd1 vccd1 hold566/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 _2907_/X vssd1 vssd1 vccd1 vccd1 _3435_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1699_ _1697_/C _1698_/Y _3462_/D vssd1 vssd1 vccd1 vccd1 _3573_/D sky130_fd_sc_hd__a21oi_1
X_3438_ _3438_/CLK _3438_/D vssd1 vssd1 vccd1 vccd1 _3438_/Q sky130_fd_sc_hd__dfxtp_1
Xhold599 _2885_/X vssd1 vssd1 vccd1 vccd1 _3415_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _3429_/CLK _3369_/D vssd1 vssd1 vccd1 vccd1 _3369_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput42 _2561_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_12
XANTENNA__2797__S _2799_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput53 _3650_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_12
Xoutput64 _2527_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_12
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_58_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2561__A _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2740_ hold37/X _2760_/B vssd1 vssd1 vccd1 vccd1 _2749_/S sky130_fd_sc_hd__or2_4
XFILLER_0_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2671_ hold241/X _2804_/A1 _2676_/S vssd1 vssd1 vccd1 vccd1 _2671_/X sky130_fd_sc_hd__mux2_1
X_1622_ _1557_/A _2576_/A _1622_/S vssd1 vssd1 vccd1 vccd1 _1622_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1624__B _1624_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3223_ _3509_/CLK _3223_/D vssd1 vssd1 vccd1 vccd1 _3223_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3154_ _3424_/CLK _3154_/D vssd1 vssd1 vccd1 vccd1 _3154_/Q sky130_fd_sc_hd__dfxtp_1
X_3085_ _3122_/A vssd1 vssd1 vccd1 vccd1 _3085_/Y sky130_fd_sc_hd__inv_2
X_2105_ _2105_/A _2105_/B vssd1 vssd1 vccd1 vccd1 _2110_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2036_ _2034_/X _2035_/X _2036_/S vssd1 vssd1 vccd1 vccd1 _2036_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2938_ _3127_/A vssd1 vssd1 vccd1 vccd1 _2938_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2869_ hold524/X _2355_/B _2870_/S vssd1 vssd1 vccd1 vccd1 _2869_/X sky130_fd_sc_hd__mux2_1
Xhold341 _3291_/Q vssd1 vssd1 vccd1 vccd1 hold341/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold330 _3295_/Q vssd1 vssd1 vccd1 vccd1 hold330/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 _2765_/X vssd1 vssd1 vccd1 vccd1 _3293_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 _2777_/X vssd1 vssd1 vccd1 vccd1 _3304_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 _3619_/Q vssd1 vssd1 vccd1 vccd1 hold396/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _3210_/Q vssd1 vssd1 vccd1 vccd1 hold374/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 _3634_/Q vssd1 vssd1 vccd1 vccd1 _1557_/A sky130_fd_sc_hd__clkbuf_2
Xhold1041 wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1030 _3349_/Q vssd1 vssd1 vccd1 vccd1 _2378_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1052 _3529_/Q vssd1 vssd1 vccd1 vccd1 hold1052/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2005__S0 _2221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2556__A _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1610__D input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2723_ _2804_/A1 hold190/X _2728_/S vssd1 vssd1 vccd1 vccd1 _2723_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_81_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2654_ _2356_/B hold586/X _2654_/S vssd1 vssd1 vccd1 vccd1 _2654_/X sky130_fd_sc_hd__mux2_1
X_2585_ hold405/X _2805_/A1 _2589_/S vssd1 vssd1 vccd1 vccd1 _2585_/X sky130_fd_sc_hd__mux2_1
X_1605_ _3054_/A vssd1 vssd1 vccd1 vccd1 _1605_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout128 _3057_/A vssd1 vssd1 vccd1 vccd1 _3061_/A sky130_fd_sc_hd__buf_4
Xfanout106 hold117/X vssd1 vssd1 vccd1 vccd1 _2804_/A1 sky130_fd_sc_hd__buf_4
Xfanout117 _3112_/A vssd1 vssd1 vccd1 vccd1 _3067_/A sky130_fd_sc_hd__clkbuf_4
X_3206_ _3330_/CLK _3206_/D vssd1 vssd1 vccd1 vccd1 _3206_/Q sky130_fd_sc_hd__dfxtp_1
X_3137_ _3332_/CLK _3137_/D vssd1 vssd1 vccd1 vccd1 _3137_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_hold1018_A _3577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3068_ _3069_/A vssd1 vssd1 vccd1 vccd1 _3068_/Y sky130_fd_sc_hd__inv_2
X_2019_ _2036_/S _2015_/X _2315_/A1 vssd1 vssd1 vccd1 vccd1 _2019_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_18_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2483__S0 _2532_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold171 _3200_/Q vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 _2744_/X vssd1 vssd1 vccd1 vccd1 _3274_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _3209_/Q vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 _2706_/X vssd1 vssd1 vccd1 vccd1 _3242_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2863__A1 _2098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2370_ _2370_/A vssd1 vssd1 vccd1 vccd1 _2370_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2529__S1 _1943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2706_ _2808_/A1 hold192/X _2707_/S vssd1 vssd1 vccd1 vccd1 _2706_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2637_ _2109_/B hold702/X _2643_/S vssd1 vssd1 vccd1 vccd1 _2637_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout118_A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2568_ hold27/A hold10/A vssd1 vssd1 vccd1 vccd1 _2568_/X sky130_fd_sc_hd__or2_1
XANTENNA__2895__S _2900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2499_ _3408_/Q _3399_/Q _3390_/Q _3435_/Q _1944_/B _1943_/A vssd1 vssd1 vccd1 vccd1
+ _2499_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_49_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2781__A0 _2801_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3429_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1870_ _1869_/X _1848_/B _1847_/A _1836_/A vssd1 vssd1 vccd1 vccd1 _1870_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_83_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2447__S0 _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3540_ _3573_/CLK _3540_/D _3034_/Y vssd1 vssd1 vccd1 vccd1 _3540_/Q sky130_fd_sc_hd__dfrtp_1
Xhold918 _3456_/Q vssd1 vssd1 vccd1 vccd1 _2270_/B sky130_fd_sc_hd__buf_1
Xhold907 _2282_/X vssd1 vssd1 vccd1 vccd1 _3457_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3471_ _3575_/CLK _3471_/D _2965_/Y vssd1 vssd1 vccd1 vccd1 _3471_/Q sky130_fd_sc_hd__dfrtp_1
Xhold929 _3439_/Q vssd1 vssd1 vccd1 vccd1 hold929/X sky130_fd_sc_hd__dlygate4sd3_1
X_2422_ _3607_/Q _2435_/A _2419_/X _2420_/X vssd1 vssd1 vccd1 vccd1 _2422_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_19_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2353_ _1571_/Y _1932_/A _1923_/A _3344_/Q vssd1 vssd1 vccd1 vccd1 _2353_/X sky130_fd_sc_hd__a211o_1
X_2284_ _2270_/B _2270_/C _2283_/Y vssd1 vssd1 vccd1 vccd1 _2284_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_79_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2827__A1 _2357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1999_ _1999_/A vssd1 vssd1 vccd1 vccd1 _1999_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2763__A0 _2803_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2818__A1 _2355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2809__A1 _2406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2564__A _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2971_ _3061_/A vssd1 vssd1 vccd1 vccd1 _2971_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_56_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1922_ _1922_/A _2613_/B _2162_/B vssd1 vssd1 vccd1 vccd1 _1924_/B sky130_fd_sc_hd__or3b_1
X_1853_ _1853_/A _1859_/A _1859_/B vssd1 vssd1 vccd1 vccd1 _1853_/X sky130_fd_sc_hd__and3_1
XFILLER_0_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1784_ _2123_/A _1784_/B _1784_/C _1784_/D vssd1 vssd1 vccd1 vccd1 _1792_/A sky130_fd_sc_hd__and4_1
XANTENNA__2745__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3523_ _3532_/CLK _3523_/D _3017_/Y vssd1 vssd1 vccd1 vccd1 _3523_/Q sky130_fd_sc_hd__dfrtp_1
Xhold737 _2886_/X vssd1 vssd1 vccd1 vccd1 _3416_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold704 _3373_/Q vssd1 vssd1 vccd1 vccd1 hold704/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 _2606_/X vssd1 vssd1 vccd1 vccd1 _3156_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 _3184_/Q vssd1 vssd1 vccd1 vccd1 hold726/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3454_ _3632_/CLK hold3/X _2948_/Y vssd1 vssd1 vccd1 vccd1 _3454_/Q sky130_fd_sc_hd__dfrtp_2
Xhold759 _2872_/X vssd1 vssd1 vccd1 vccd1 _3403_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold748 _3160_/Q vssd1 vssd1 vccd1 vccd1 hold748/X sky130_fd_sc_hd__dlygate4sd3_1
X_2405_ hold45/X hold98/X hold95/X vssd1 vssd1 vccd1 vccd1 _3587_/D sky130_fd_sc_hd__and3_1
X_3385_ _3438_/CLK _3385_/D vssd1 vssd1 vccd1 vccd1 _3385_/Q sky130_fd_sc_hd__dfxtp_1
X_2336_ _2336_/A _2336_/B vssd1 vssd1 vccd1 vccd1 _2336_/Y sky130_fd_sc_hd__nor2_1
X_2267_ _2263_/X _2267_/B _2267_/C _2267_/D vssd1 vssd1 vccd1 vccd1 _2267_/X sky130_fd_sc_hd__and4b_1
XFILLER_0_1_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2198_ hold36/X _2198_/B vssd1 vssd1 vccd1 vccd1 _2205_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_62_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout98_A _3483_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__clkbuf_4
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__clkbuf_4
Xhold97 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2727__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _3434_/CLK _3170_/D vssd1 vssd1 vccd1 vccd1 _3170_/Q sky130_fd_sc_hd__dfxtp_1
X_2121_ _2121_/A _3496_/Q vssd1 vssd1 vccd1 vccd1 _2123_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_83_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2052_ _2315_/A1 _2050_/X _2051_/Y _2046_/Y vssd1 vssd1 vccd1 vccd1 _2319_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_29_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2954_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2954_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2885_ _2101_/Y hold598/X _2890_/S vssd1 vssd1 vccd1 vccd1 _2885_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1905_ _1924_/A _1905_/B _1905_/C vssd1 vssd1 vccd1 vccd1 _3519_/D sky130_fd_sc_hd__and3_1
XANTENNA__2718__A0 _2406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1836_ _1836_/A _2228_/B vssd1 vssd1 vccd1 vccd1 _1837_/A sky130_fd_sc_hd__nor2_4
Xhold501 _2827_/X vssd1 vssd1 vccd1 vccd1 _3359_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1767_ hold778/X hold846/X _1767_/S vssd1 vssd1 vccd1 vccd1 _1767_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2194__A1 _2219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold523 _2838_/X vssd1 vssd1 vccd1 vccd1 _3369_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 _3426_/Q vssd1 vssd1 vccd1 vccd1 hold512/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 _2816_/X vssd1 vssd1 vccd1 vccd1 _3339_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 _3400_/Q vssd1 vssd1 vccd1 vccd1 hold534/X sky130_fd_sc_hd__dlygate4sd3_1
X_3506_ _3509_/CLK _3506_/D _3000_/Y vssd1 vssd1 vccd1 vccd1 _3506_/Q sky130_fd_sc_hd__dfrtp_1
Xhold567 _2889_/X vssd1 vssd1 vccd1 vccd1 _3419_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 _3189_/Q vssd1 vssd1 vccd1 vccd1 hold578/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 _3358_/Q vssd1 vssd1 vccd1 vccd1 hold556/X sky130_fd_sc_hd__dlygate4sd3_1
X_1698_ _1698_/A _1698_/B vssd1 vssd1 vccd1 vccd1 _1698_/Y sky130_fd_sc_hd__nand2_1
X_3437_ _3521_/CLK _3437_/D vssd1 vssd1 vccd1 vccd1 _3437_/Q sky130_fd_sc_hd__dfxtp_1
Xhold589 _2813_/X vssd1 vssd1 vccd1 vccd1 _3336_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _3619_/CLK _3368_/D vssd1 vssd1 vccd1 vccd1 _3368_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2319_ _2319_/A _2319_/B vssd1 vssd1 vccd1 vccd1 _2321_/A sky130_fd_sc_hd__nor2_1
X_3299_ _3319_/CLK _3299_/D vssd1 vssd1 vccd1 vccd1 _3299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1982__S _2036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput43 _2564_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_12
Xoutput54 _3651_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_12
Xoutput65 _2540_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_12
XFILLER_0_85_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2670_ hold374/X _2803_/A1 _2676_/S vssd1 vssd1 vccd1 vccd1 _2670_/X sky130_fd_sc_hd__mux2_1
X_1621_ _1950_/A _2399_/A _1622_/S vssd1 vssd1 vccd1 vccd1 _1621_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3222_ _3330_/CLK _3222_/D vssd1 vssd1 vccd1 vccd1 _3222_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3153_ _3555_/CLK _3153_/D _2917_/Y vssd1 vssd1 vccd1 vccd1 _3153_/Q sky130_fd_sc_hd__dfrtp_1
X_2104_ _2383_/B _2104_/B vssd1 vssd1 vccd1 vccd1 _2105_/B sky130_fd_sc_hd__xor2_1
X_3084_ _3090_/A vssd1 vssd1 vccd1 vccd1 _3084_/Y sky130_fd_sc_hd__inv_2
X_2035_ hold163/X hold182/X hold171/X hold174/X _2045_/S0 _2045_/S1 vssd1 vssd1 vccd1
+ vccd1 _2035_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2100__B2 _2064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2937_ _3127_/A vssd1 vssd1 vccd1 vccd1 _2937_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2898__S _2900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2868_ hold534/X _2357_/B _2870_/S vssd1 vssd1 vccd1 vccd1 _2868_/X sky130_fd_sc_hd__mux2_1
X_2799_ hold47/X hold30/X _2799_/S vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__mux2_1
XFILLER_0_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold320 _2675_/X vssd1 vssd1 vccd1 vccd1 _3215_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1819_ _3551_/Q _1809_/B _1824_/A _1742_/B vssd1 vssd1 vccd1 vccd1 _1819_/X sky130_fd_sc_hd__o211a_1
Xhold342 _2763_/X vssd1 vssd1 vccd1 vccd1 _3291_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 _2767_/X vssd1 vssd1 vccd1 vccd1 _3295_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 _3132_/Q vssd1 vssd1 vccd1 vccd1 hold353/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold386 _3257_/Q vssd1 vssd1 vccd1 vccd1 hold386/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 _2670_/X vssd1 vssd1 vccd1 vccd1 _3210_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 _1622_/X vssd1 vssd1 vccd1 vccd1 _3634_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold397 _3230_/Q vssd1 vssd1 vccd1 vccd1 hold397/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 input13/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1020 _1716_/Y vssd1 vssd1 vccd1 vccd1 _1728_/D1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1053 _3472_/Q vssd1 vssd1 vccd1 vccd1 hold943/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1669__A0 _2401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2005__S1 _2219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2722_ _2803_/A1 hold321/X _2728_/S vssd1 vssd1 vccd1 vccd1 _2722_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2653_ _2355_/B hold580/X _2654_/S vssd1 vssd1 vccd1 vccd1 _2653_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2584_ hold214/X _2804_/A1 _2589_/S vssd1 vssd1 vccd1 vccd1 _2584_/X sky130_fd_sc_hd__mux2_1
X_1604_ _1809_/A vssd1 vssd1 vccd1 vccd1 _1816_/B sky130_fd_sc_hd__inv_2
Xfanout129 input2/X vssd1 vssd1 vccd1 vccd1 _3057_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout107 hold117/X vssd1 vssd1 vccd1 vccd1 _2401_/A sky130_fd_sc_hd__clkbuf_4
Xfanout118 _3112_/A vssd1 vssd1 vccd1 vccd1 _3129_/A sky130_fd_sc_hd__buf_8
X_3205_ _3509_/CLK _3205_/D vssd1 vssd1 vccd1 vccd1 _3205_/Q sky130_fd_sc_hd__dfxtp_1
X_3136_ _3509_/CLK _3136_/D vssd1 vssd1 vccd1 vccd1 _3136_/Q sky130_fd_sc_hd__dfxtp_1
X_3067_ _3067_/A vssd1 vssd1 vccd1 vccd1 _3067_/Y sky130_fd_sc_hd__inv_2
X_2018_ _2017_/X _2016_/X _2036_/S vssd1 vssd1 vccd1 vccd1 _2018_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2483__S1 _2532_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold150 input5/X vssd1 vssd1 vccd1 vccd1 _1657_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 _3301_/Q vssd1 vssd1 vccd1 vccd1 hold161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 _3238_/Q vssd1 vssd1 vccd1 vccd1 hold194/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _2659_/X vssd1 vssd1 vccd1 vccd1 _3200_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _2669_/X vssd1 vssd1 vccd1 vccd1 _3209_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold477_A _3517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output61_A _2487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2567__A _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2303__A1 _2400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3319_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2705_ _2807_/A1 hold421/X _2707_/S vssd1 vssd1 vccd1 vccd1 _2705_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2636_ _2098_/S hold746/X _2643_/S vssd1 vssd1 vccd1 vccd1 _2636_/X sky130_fd_sc_hd__mux2_1
X_2567_ _2574_/A _2567_/B vssd1 vssd1 vccd1 vccd1 _2567_/X sky130_fd_sc_hd__and2_2
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2498_ _1908_/D _2497_/X _2492_/X vssd1 vssd1 vccd1 vccd1 _2498_/X sky130_fd_sc_hd__a21o_1
X_3119_ _3122_/A vssd1 vssd1 vccd1 vccd1 _3119_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1990__S _2055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2447__S1 _1943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2772__A1 _2802_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold919 _2284_/X vssd1 vssd1 vccd1 vccd1 _3456_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold908 _3574_/Q vssd1 vssd1 vccd1 vccd1 hold908/X sky130_fd_sc_hd__dlygate4sd3_1
X_3470_ _3574_/CLK _3470_/D _2964_/Y vssd1 vssd1 vccd1 vccd1 _3470_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2421_ _2421_/A _2421_/B vssd1 vssd1 vccd1 vccd1 _2507_/C sky130_fd_sc_hd__nand2_2
X_2352_ _1571_/Y _1932_/A _3513_/Q _1572_/Y _2351_/X vssd1 vssd1 vccd1 vccd1 _2352_/X
+ sky130_fd_sc_hd__o221a_1
X_2283_ _2283_/A _2283_/B vssd1 vssd1 vccd1 vccd1 _2283_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1998_ _2315_/A1 _1993_/X _1997_/X vssd1 vssd1 vccd1 vccd1 _1999_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_70_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3599_ _3600_/CLK _3599_/D _3090_/Y vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__dfrtp_1
X_2619_ _2104_/B hold760/X _2623_/S vssd1 vssd1 vccd1 vccd1 _2619_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_65_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1985__S _2036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2754__A1 _2804_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2970_ _3061_/A vssd1 vssd1 vccd1 vccd1 _2970_/Y sky130_fd_sc_hd__inv_2
X_1921_ _1918_/B _1911_/Y _1918_/X vssd1 vssd1 vccd1 vccd1 _3515_/D sky130_fd_sc_hd__o21ba_1
XFILLER_0_29_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1852_ _1859_/A _1859_/B vssd1 vssd1 vccd1 vccd1 _1852_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1908__B _3577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1783_ _3553_/Q _2122_/B vssd1 vssd1 vccd1 vccd1 _1784_/D sky130_fd_sc_hd__xor2_1
XFILLER_0_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold705 _2843_/X vssd1 vssd1 vccd1 vccd1 _3373_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 _2638_/X vssd1 vssd1 vccd1 vccd1 _3184_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold716 _3431_/Q vssd1 vssd1 vccd1 vccd1 hold716/X sky130_fd_sc_hd__dlygate4sd3_1
X_3522_ _3602_/CLK _3522_/D _3016_/Y vssd1 vssd1 vccd1 vccd1 _3522_/Q sky130_fd_sc_hd__dfrtp_4
X_3453_ _3632_/CLK hold26/X _2947_/Y vssd1 vssd1 vccd1 vccd1 _3453_/Q sky130_fd_sc_hd__dfrtp_1
Xhold738 _3389_/Q vssd1 vssd1 vccd1 vccd1 hold738/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 _2610_/X vssd1 vssd1 vccd1 vccd1 _3160_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2404_ hold87/X hold98/X hold95/X vssd1 vssd1 vccd1 vccd1 _3586_/D sky130_fd_sc_hd__and3_1
X_3384_ _3607_/CLK _3384_/D _2932_/Y vssd1 vssd1 vccd1 vccd1 _3384_/Q sky130_fd_sc_hd__dfrtp_1
X_2335_ _2335_/A1 _2363_/A _3381_/Q vssd1 vssd1 vccd1 vccd1 _2336_/B sky130_fd_sc_hd__a21oi_1
X_2266_ _3630_/Q _1594_/Y _2270_/B _2550_/A _2261_/Y vssd1 vssd1 vccd1 vccd1 _2267_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2197_ hold36/X _2198_/B vssd1 vssd1 vccd1 vccd1 _2208_/B sky130_fd_sc_hd__and2_2
XANTENNA__2681__A0 _2803_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2736__A1 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold32 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 input8/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__clkbuf_4
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__clkbuf_4
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__buf_2
XFILLER_0_85_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2604__S _2612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3532_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2120_ _2121_/A _3496_/Q vssd1 vssd1 vccd1 vccd1 _2123_/B sky130_fd_sc_hd__or2_1
XANTENNA__2575__A _2576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2051_ _2036_/S _2047_/X _2315_/A1 vssd1 vssd1 vccd1 vccd1 _2051_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__2663__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2953_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2953_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1904_ _1904_/A _2613_/B vssd1 vssd1 vccd1 vccd1 _1905_/C sky130_fd_sc_hd__or2_1
X_2884_ _2108_/Y hold596/X _2890_/S vssd1 vssd1 vccd1 vccd1 _2884_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1835_ _3540_/Q hold813/X _1835_/S vssd1 vssd1 vccd1 vccd1 _1835_/X sky130_fd_sc_hd__mux2_1
Xhold502 _3394_/Q vssd1 vssd1 vccd1 vccd1 hold502/X sky130_fd_sc_hd__dlygate4sd3_1
X_1766_ hold957/X _1743_/Y _1765_/X vssd1 vssd1 vccd1 vccd1 _1766_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2194__A2 _2221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold513 _2897_/X vssd1 vssd1 vccd1 vccd1 _3426_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 _3401_/Q vssd1 vssd1 vccd1 vccd1 hold524/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold535 _2868_/X vssd1 vssd1 vccd1 vccd1 _3400_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3505_ _3509_/CLK _3505_/D _2999_/Y vssd1 vssd1 vccd1 vccd1 _3505_/Q sky130_fd_sc_hd__dfrtp_1
Xhold579 _2643_/X vssd1 vssd1 vccd1 vccd1 _3189_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 _3143_/Q vssd1 vssd1 vccd1 vccd1 hold568/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 _3377_/Q vssd1 vssd1 vccd1 vccd1 hold546/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 _2826_/X vssd1 vssd1 vccd1 vccd1 _3358_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1697_ _1697_/A _1697_/B _1697_/C vssd1 vssd1 vccd1 vccd1 _1697_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3436_ _3521_/CLK _3436_/D vssd1 vssd1 vccd1 vccd1 _3436_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _3516_/CLK _3367_/D vssd1 vssd1 vccd1 vccd1 _3367_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ _2316_/A _2316_/B _2316_/Y _2317_/X vssd1 vssd1 vccd1 vccd1 _2322_/A sky130_fd_sc_hd__o211ai_1
X_3298_ _3318_/CLK _3298_/D vssd1 vssd1 vccd1 vccd1 _3298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2249_ _2249_/A _3464_/Q _3463_/Q _2249_/D vssd1 vssd1 vccd1 vccd1 _2249_/X sky130_fd_sc_hd__or4_1
XANTENNA__2654__A0 _2356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput55 _3652_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_12
Xoutput66 _2552_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_12
Xoutput44 _2567_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_12
XFILLER_0_37_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1620__A1 _2400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1620_ _1888_/A _2400_/A _1622_/S vssd1 vssd1 vccd1 vccd1 _1620_/X sky130_fd_sc_hd__mux2_1
X_3221_ _3329_/CLK _3221_/D vssd1 vssd1 vccd1 vccd1 _3221_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1687__A1 _2576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3152_ _3550_/CLK _3152_/D _2916_/Y vssd1 vssd1 vccd1 vccd1 _3152_/Q sky130_fd_sc_hd__dfrtp_1
X_2103_ _2065_/Y _2090_/B _2102_/X _2067_/B vssd1 vssd1 vccd1 vccd1 _2103_/Y sky130_fd_sc_hd__a211oi_4
X_3083_ _3122_/A vssd1 vssd1 vccd1 vccd1 _3083_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2636__A0 _2098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2034_ hold179/X hold186/X hold176/X hold184/X _2045_/S0 _2045_/S1 vssd1 vssd1 vccd1
+ vccd1 _2034_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2936_ _3127_/A vssd1 vssd1 vccd1 vccd1 _2936_/Y sky130_fd_sc_hd__inv_2
X_2867_ hold506/X _2360_/B _2870_/S vssd1 vssd1 vccd1 vccd1 _2867_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1818_ _1818_/A _1818_/B vssd1 vssd1 vccd1 vccd1 _1824_/A sky130_fd_sc_hd__and2_1
X_2798_ hold251/X _2808_/A1 _2799_/S vssd1 vssd1 vccd1 vccd1 _2798_/X sky130_fd_sc_hd__mux2_1
Xhold310 _2737_/X vssd1 vssd1 vccd1 vccd1 _3268_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 _3270_/Q vssd1 vssd1 vccd1 vccd1 hold343/X sky130_fd_sc_hd__dlygate4sd3_1
X_1749_ _1811_/S _1749_/B _1769_/B vssd1 vssd1 vccd1 vccd1 _1749_/X sky130_fd_sc_hd__or3_1
XFILLER_0_7_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold321 _3255_/Q vssd1 vssd1 vccd1 vccd1 hold321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 _3320_/Q vssd1 vssd1 vccd1 vccd1 hold332/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 _2724_/X vssd1 vssd1 vccd1 vccd1 _3257_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 _3258_/Q vssd1 vssd1 vccd1 vccd1 hold376/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 _3609_/Q vssd1 vssd1 vccd1 vccd1 _1572_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 _2583_/X vssd1 vssd1 vccd1 vccd1 _3132_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3419_ _3429_/CLK _3419_/D vssd1 vssd1 vccd1 vccd1 _3419_/Q sky130_fd_sc_hd__dfxtp_1
Xhold398 _2693_/X vssd1 vssd1 vccd1 vccd1 _3230_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1678__A1 hold59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2875__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1021 _3449_/Q vssd1 vssd1 vccd1 vccd1 _1717_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1010 _1800_/X vssd1 vssd1 vccd1 vccd1 _1801_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 _1612_/X vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1054 _3492_/Q vssd1 vssd1 vccd1 vccd1 hold985/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 _3602_/Q vssd1 vssd1 vccd1 vccd1 hold466/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3104__A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2627__A0 _2109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1993__S _2036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2618__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2572__B hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2721_ _2802_/A1 hold179/X _2728_/S vssd1 vssd1 vccd1 vccd1 _2721_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2652_ _2357_/B hold504/X _2654_/S vssd1 vssd1 vccd1 vccd1 _2652_/X sky130_fd_sc_hd__mux2_1
X_2583_ hold353/X _2803_/A1 _2589_/S vssd1 vssd1 vccd1 vccd1 _2583_/X sky130_fd_sc_hd__mux2_1
X_1603_ _2211_/A vssd1 vssd1 vccd1 vccd1 _2177_/A sky130_fd_sc_hd__inv_2
XFILLER_0_22_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout108 hold120/X vssd1 vssd1 vccd1 vccd1 _2803_/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_10_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout119 _3112_/A vssd1 vssd1 vccd1 vccd1 _3049_/A sky130_fd_sc_hd__buf_6
XFILLER_0_10_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3204_ _3329_/CLK _3204_/D vssd1 vssd1 vccd1 vccd1 _3204_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2857__A0 _2360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3135_ _3329_/CLK _3135_/D vssd1 vssd1 vccd1 vccd1 _3135_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2609__A0 _2360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3066_ _3067_/A vssd1 vssd1 vccd1 vccd1 _3066_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2017_ _3247_/Q _3319_/Q _3310_/Q _3301_/Q _2221_/B _2219_/A vssd1 vssd1 vccd1 vccd1
+ _2017_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_64_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2919_ _3101_/A vssd1 vssd1 vccd1 vccd1 _2919_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2388__A2 _1769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2702__S _2707_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold151 _1674_/B vssd1 vssd1 vccd1 vccd1 _1659_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 _3281_/Q vssd1 vssd1 vccd1 vccd1 hold140/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 _2774_/X vssd1 vssd1 vccd1 vccd1 _3301_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _2702_/X vssd1 vssd1 vccd1 vccd1 _3238_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _3227_/Q vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 hold173/A vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__buf_1
XANTENNA__1994__S1 _2195_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2848__A0 _2355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2612__S _2612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2839__A0 _2356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2704_ _2806_/A1 hold392/X _2707_/S vssd1 vssd1 vccd1 vccd1 _2704_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2635_ _2358_/B hold708/X _2643_/S vssd1 vssd1 vccd1 vccd1 _2635_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2566_ _3452_/Q _2510_/B _2559_/X _2565_/X vssd1 vssd1 vccd1 vccd1 _2567_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_10_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2497_ _2495_/X _2496_/X _2493_/X _2494_/X _3517_/Q _3518_/Q vssd1 vssd1 vccd1 vccd1
+ _2497_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3118_ _3129_/A vssd1 vssd1 vccd1 vccd1 _3118_/Y sky130_fd_sc_hd__inv_2
XANTENNA_hold1023_A _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3049_ _3049_/A vssd1 vssd1 vccd1 vccd1 _3049_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_81_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2432__S _2546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2297__A1 _2406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2607__S _2612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_48_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3434_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout90 hold914/X vssd1 vssd1 vccd1 vccd1 _2225_/A sky130_fd_sc_hd__buf_2
XFILLER_0_24_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold909 _3485_/Q vssd1 vssd1 vccd1 vccd1 hold909/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2420_ _2421_/A _2421_/B vssd1 vssd1 vccd1 vccd1 _2420_/X sky130_fd_sc_hd__and2_1
XFILLER_0_19_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2351_ _1574_/Y _1941_/S _2349_/X _2350_/X vssd1 vssd1 vccd1 vccd1 _2351_/X sky130_fd_sc_hd__a31o_1
X_2282_ _2270_/A _2283_/B _2281_/Y vssd1 vssd1 vccd1 vccd1 _2282_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2517__S _2546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1997_ _2225_/A _1997_/B vssd1 vssd1 vccd1 vccd1 _1997_/X sky130_fd_sc_hd__and2b_1
XANTENNA_fanout123_A _3124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1657__A _1657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2618_ _2105_/A hold620/X _2623_/S vssd1 vssd1 vccd1 vccd1 _2618_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3598_ _3600_/CLK hold88/X _3089_/Y vssd1 vssd1 vccd1 vccd1 _3598_/Q sky130_fd_sc_hd__dfrtp_1
X_2549_ _3588_/Q hold95/A _2410_/X _3382_/Q _2548_/X vssd1 vssd1 vccd1 vccd1 _2549_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3112__A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2951__A _3124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2398__A _2576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2690__A1 _2802_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1920_ _1912_/B _1918_/X hold467/X _1911_/B vssd1 vssd1 vccd1 vccd1 _1920_/X sky130_fd_sc_hd__o22a_1
X_1851_ _1851_/A _1851_/B vssd1 vssd1 vccd1 vccd1 _1859_/B sky130_fd_sc_hd__and2_1
XFILLER_0_21_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3521_ _3521_/CLK _3521_/D _3015_/Y vssd1 vssd1 vccd1 vccd1 _3521_/Q sky130_fd_sc_hd__dfrtp_4
X_1782_ _2070_/A _2092_/A vssd1 vssd1 vccd1 vccd1 _2122_/B sky130_fd_sc_hd__xor2_2
Xhold717 _2903_/X vssd1 vssd1 vccd1 vccd1 _3431_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold728 _3375_/Q vssd1 vssd1 vccd1 vccd1 hold728/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold706 _3175_/Q vssd1 vssd1 vccd1 vccd1 hold706/X sky130_fd_sc_hd__dlygate4sd3_1
X_3452_ _3632_/CLK hold23/X _2946_/Y vssd1 vssd1 vccd1 vccd1 _3452_/Q sky130_fd_sc_hd__dfrtp_1
Xhold739 _2856_/X vssd1 vssd1 vccd1 vccd1 _3389_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3383_ _3589_/CLK _3383_/D _2931_/Y vssd1 vssd1 vccd1 vccd1 _3383_/Q sky130_fd_sc_hd__dfrtp_1
X_2403_ hold70/X hold98/X hold95/X vssd1 vssd1 vccd1 vccd1 _3585_/D sky130_fd_sc_hd__and3_1
X_2334_ _2334_/A _2334_/B vssd1 vssd1 vccd1 vccd1 _2334_/Y sky130_fd_sc_hd__nor2_1
X_2265_ hold80/X _1593_/Y _2271_/B _1559_/Y _2264_/X vssd1 vssd1 vccd1 vccd1 _2267_/B
+ sky130_fd_sc_hd__o221a_1
X_2196_ _2193_/A _2186_/X hold890/X vssd1 vssd1 vccd1 vccd1 _2196_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2490__B hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2710__S _2718_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3107__A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__buf_4
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 input8/X vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2672__A1 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2035__S0 _2045_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2050_ _2049_/X _2048_/X _2222_/A vssd1 vssd1 vccd1 vccd1 _2050_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2952_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2952_/Y sky130_fd_sc_hd__inv_2
X_1903_ _1901_/Y hold809/X _1935_/A vssd1 vssd1 vccd1 vccd1 _1903_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2883_ _2087_/Y hold550/X _2890_/S vssd1 vssd1 vccd1 vccd1 _2883_/X sky130_fd_sc_hd__mux2_1
X_1834_ hold827/X _3540_/Q _1835_/S vssd1 vssd1 vccd1 vccd1 _1834_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1765_ _1811_/S _3556_/Q _1769_/B vssd1 vssd1 vccd1 vccd1 _1765_/X sky130_fd_sc_hd__or3_1
XANTENNA__2530__S _2546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold514 _3396_/Q vssd1 vssd1 vccd1 vccd1 hold514/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold503 _2862_/X vssd1 vssd1 vccd1 vccd1 _3394_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 _3338_/Q vssd1 vssd1 vccd1 vccd1 hold536/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 _2869_/X vssd1 vssd1 vccd1 vccd1 _3401_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3504_ _3504_/CLK _3504_/D _2998_/Y vssd1 vssd1 vccd1 vccd1 _3504_/Q sky130_fd_sc_hd__dfrtp_1
Xhold569 _2597_/X vssd1 vssd1 vccd1 vccd1 _3143_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 _3368_/Q vssd1 vssd1 vccd1 vccd1 hold558/X sky130_fd_sc_hd__dlygate4sd3_1
X_3435_ _3438_/CLK _3435_/D vssd1 vssd1 vccd1 vccd1 _3435_/Q sky130_fd_sc_hd__dfxtp_1
X_1696_ _1697_/B _1697_/C _1695_/X vssd1 vssd1 vccd1 vccd1 _3574_/D sky130_fd_sc_hd__a21bo_1
Xhold547 _2847_/X vssd1 vssd1 vccd1 vccd1 _3377_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2026__S0 _2045_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3366_ _3431_/CLK _3366_/D vssd1 vssd1 vccd1 vccd1 _3366_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3297_ _3484_/CLK hold31/X vssd1 vssd1 vccd1 vccd1 _3297_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ _2070_/A _2121_/A _1774_/X vssd1 vssd1 vccd1 vccd1 _2317_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_57_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2248_ _2248_/A _3469_/Q _3468_/Q _3467_/Q vssd1 vssd1 vccd1 vccd1 _2249_/D sky130_fd_sc_hd__or4_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2179_ _2677_/B hold36/X _2178_/Y vssd1 vssd1 vccd1 vccd1 _2179_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2705__S _2707_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput67 _2556_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_12
Xoutput56 _3653_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_12
Xoutput45 _2570_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_12
XANTENNA__2017__S0 _2221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3220_ _3509_/CLK _3220_/D vssd1 vssd1 vccd1 vccd1 _3220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3151_ _3559_/CLK _3151_/D _2915_/Y vssd1 vssd1 vccd1 vccd1 _3151_/Q sky130_fd_sc_hd__dfrtp_1
X_2102_ _2070_/A _2096_/B _2090_/A vssd1 vssd1 vccd1 vccd1 _2102_/X sky130_fd_sc_hd__o21a_1
X_3082_ _3097_/A vssd1 vssd1 vccd1 vccd1 _3082_/Y sky130_fd_sc_hd__inv_2
X_2033_ hold792/X _2032_/Y _2055_/S vssd1 vssd1 vccd1 vccd1 _2033_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2935_ _3127_/A vssd1 vssd1 vccd1 vccd1 _2935_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2495__S0 _1918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2866_ hold718/X _2104_/B _2870_/S vssd1 vssd1 vccd1 vccd1 _2866_/X sky130_fd_sc_hd__mux2_1
X_1817_ _1886_/A _1814_/Y _1815_/X _1816_/Y vssd1 vssd1 vccd1 vccd1 _1817_/X sky130_fd_sc_hd__o22a_1
X_2797_ hold380/X _2807_/A1 _2799_/S vssd1 vssd1 vccd1 vccd1 _2797_/X sky130_fd_sc_hd__mux2_1
Xhold311 _3620_/Q vssd1 vssd1 vccd1 vccd1 hold311/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold300 _2686_/X vssd1 vssd1 vccd1 vccd1 _3224_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 _2739_/X vssd1 vssd1 vccd1 vccd1 _3270_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1748_ hold971/X _2387_/C _1747_/X vssd1 vssd1 vccd1 vccd1 _1748_/X sky130_fd_sc_hd__o21a_1
Xhold322 _2722_/X vssd1 vssd1 vccd1 vccd1 _3255_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 _2795_/X vssd1 vssd1 vccd1 vccd1 _3320_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 _3286_/Q vssd1 vssd1 vccd1 vccd1 hold366/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 _2725_/X vssd1 vssd1 vccd1 vccd1 _3258_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 _3201_/Q vssd1 vssd1 vccd1 vccd1 hold355/X sky130_fd_sc_hd__dlygate4sd3_1
X_1679_ hold390/X _2406_/A hold65/X vssd1 vssd1 vccd1 vccd1 _3600_/D sky130_fd_sc_hd__mux2_1
X_3418_ _3575_/CLK _3418_/D vssd1 vssd1 vccd1 vccd1 _3418_/Q sky130_fd_sc_hd__dfxtp_1
Xhold399 _3207_/Q vssd1 vssd1 vccd1 vccd1 hold399/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 _3239_/Q vssd1 vssd1 vccd1 vccd1 hold388/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1000 _3473_/Q vssd1 vssd1 vccd1 vccd1 _2228_/C sky130_fd_sc_hd__dlygate4sd3_1
X_3349_ _3635_/CLK _3349_/D _2924_/Y vssd1 vssd1 vccd1 vccd1 _3349_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1022 _1950_/B vssd1 vssd1 vccd1 vccd1 _1888_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1011 _1801_/X vssd1 vssd1 vccd1 vccd1 _3554_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 _2165_/B vssd1 vssd1 vccd1 vccd1 _1661_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1055 _3534_/Q vssd1 vssd1 vccd1 vccd1 hold1055/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 _3624_/Q vssd1 vssd1 vccd1 vccd1 hold102/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold150_A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2866__A1 _2104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2720_ _2801_/A1 hold255/X _2728_/S vssd1 vssd1 vccd1 vccd1 _2720_/X sky130_fd_sc_hd__mux2_1
X_2651_ _2360_/B hold660/X _2654_/S vssd1 vssd1 vccd1 vccd1 _2651_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1602_ _1935_/A vssd1 vssd1 vccd1 vccd1 _1924_/A sky130_fd_sc_hd__inv_2
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2582_ hold186/X _2802_/A1 _2589_/S vssd1 vssd1 vccd1 vccd1 _2582_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout109 hold120/X vssd1 vssd1 vccd1 vccd1 _2400_/A sky130_fd_sc_hd__clkbuf_4
X_3203_ _3329_/CLK _3203_/D vssd1 vssd1 vccd1 vccd1 _3203_/Q sky130_fd_sc_hd__dfxtp_1
X_3134_ _3326_/CLK _3134_/D vssd1 vssd1 vccd1 vccd1 _3134_/Q sky130_fd_sc_hd__dfxtp_1
X_3065_ _3067_/A vssd1 vssd1 vccd1 vccd1 _3065_/Y sky130_fd_sc_hd__inv_2
X_2016_ hold155/X hold165/X hold159/X hold167/X _2221_/B _2219_/A vssd1 vssd1 vccd1
+ vccd1 _2016_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_70_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2918_ _3090_/A vssd1 vssd1 vccd1 vccd1 _2918_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2849_ _2356_/B hold590/X _2849_/S vssd1 vssd1 vccd1 vccd1 _2849_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold130 _2782_/X vssd1 vssd1 vccd1 vccd1 _3308_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold152 _2421_/A vssd1 vssd1 vccd1 vccd1 _2416_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 _2752_/X vssd1 vssd1 vccd1 vccd1 _3281_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _2690_/X vssd1 vssd1 vccd1 vccd1 _3227_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 _3218_/Q vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 _3326_/Q vssd1 vssd1 vccd1 vccd1 hold174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 _3260_/Q vssd1 vssd1 vccd1 vccd1 hold196/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2954__A _3124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2784__A0 _2804_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2703_ _2805_/A1 hold388/X _2707_/S vssd1 vssd1 vccd1 vccd1 _2703_/X sky130_fd_sc_hd__mux2_1
X_2634_ _3520_/Q _3519_/Q _2871_/C _2810_/B vssd1 vssd1 vccd1 vccd1 _2643_/S sky130_fd_sc_hd__or4b_4
XANTENNA__2104__A _2383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2565_ _3632_/Q hold10/A vssd1 vssd1 vccd1 vccd1 _2565_/X sky130_fd_sc_hd__or2_1
XFILLER_0_2_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1943__A _1943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2496_ _3375_/Q _3357_/Q _3366_/Q _3194_/Q _1918_/B _1912_/B vssd1 vssd1 vccd1 vccd1
+ _2496_/X sky130_fd_sc_hd__mux4_1
X_3117_ _3129_/A vssd1 vssd1 vccd1 vccd1 _3117_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3048_ _3049_/A vssd1 vssd1 vccd1 vccd1 _3048_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_65_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2713__S _2718_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2766__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout91 _3485_/Q vssd1 vssd1 vccd1 vccd1 _2036_/S sky130_fd_sc_hd__clkbuf_8
Xfanout80 _2121_/A vssd1 vssd1 vccd1 vccd1 _2092_/A sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_17_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3590_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2350_ _1572_/Y _3513_/Q _2349_/B _2349_/A vssd1 vssd1 vccd1 vccd1 _2350_/X sky130_fd_sc_hd__a22o_1
X_2281_ _2283_/A _2281_/B vssd1 vssd1 vccd1 vccd1 _2281_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2445__C1 _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2460__A2 hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2748__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1996_ _1995_/X _1994_/X _2222_/A vssd1 vssd1 vccd1 vccd1 _1997_/B sky130_fd_sc_hd__mux2_1
XANTENNA__2533__S _3517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1657__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout116_A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2617_ _2109_/B hold762/X _2623_/S vssd1 vssd1 vccd1 vccd1 _2617_/X sky130_fd_sc_hd__mux2_1
X_3597_ _3600_/CLK _3597_/D _3088_/Y vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__dfrtp_1
X_2548_ _3382_/Q _1675_/X _2409_/Y _3600_/Q vssd1 vssd1 vccd1 vccd1 _2548_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2479_ _3443_/Q hold21/A _2478_/X _2574_/A vssd1 vssd1 vccd1 vccd1 _2479_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_33_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1850_ _1850_/A _1865_/A _1865_/B vssd1 vssd1 vccd1 vccd1 _1851_/B sky130_fd_sc_hd__and3_1
XFILLER_0_4_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1781_ _2092_/A _3552_/Q vssd1 vssd1 vccd1 vccd1 _1784_/C sky130_fd_sc_hd__nand2_1
X_3520_ _3521_/CLK _3520_/D _3014_/Y vssd1 vssd1 vccd1 vccd1 _3520_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_24_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1908__D _1908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold718 _3398_/Q vssd1 vssd1 vccd1 vccd1 hold718/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold707 _2628_/X vssd1 vssd1 vccd1 vccd1 _3175_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3451_ _3633_/CLK hold79/X _2945_/Y vssd1 vssd1 vccd1 vccd1 _3451_/Q sky130_fd_sc_hd__dfrtp_1
Xhold729 _2845_/X vssd1 vssd1 vccd1 vccd1 _3375_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3382_ _3607_/CLK _3382_/D _2930_/Y vssd1 vssd1 vccd1 vccd1 _3382_/Q sky130_fd_sc_hd__dfrtp_1
X_2402_ hold75/X hold98/X hold95/X vssd1 vssd1 vccd1 vccd1 _3584_/D sky130_fd_sc_hd__and3_1
XANTENNA__2902__A0 _2358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2333_ _1923_/A _2363_/A _3382_/Q vssd1 vssd1 vccd1 vccd1 _2334_/B sky130_fd_sc_hd__a21oi_1
X_2264_ _2550_/A _3456_/Q hold806/X _1558_/Y vssd1 vssd1 vccd1 vccd1 _2264_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2195_ _2195_/A1 _2193_/Y _2194_/Y _2227_/A vssd1 vssd1 vccd1 vccd1 _2195_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_46_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1979_ hold788/X _1978_/X _2055_/S vssd1 vssd1 vccd1 vccd1 _1979_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3649_ _3655_/A vssd1 vssd1 vccd1 vccd1 _3649_/X sky130_fd_sc_hd__buf_1
XFILLER_0_87_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__clkbuf_8
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__clkbuf_4
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3123__A _3124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2424__A2 hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2035__S1 _2045_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2951_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2951_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1902_ _1902_/A _1905_/B vssd1 vssd1 vccd1 vccd1 _1902_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_32_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3622_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2882_ _2097_/X hold744/X _2890_/S vssd1 vssd1 vccd1 vccd1 _2882_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1833_ hold844/X hold827/X _1833_/S vssd1 vssd1 vccd1 vccd1 _3541_/D sky130_fd_sc_hd__mux2_1
X_1764_ _1761_/B _2387_/C _1763_/X vssd1 vssd1 vccd1 vccd1 _1764_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_52_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold515 _2864_/X vssd1 vssd1 vccd1 vccd1 _3396_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold526 _3428_/Q vssd1 vssd1 vccd1 vccd1 hold526/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold504 _3196_/Q vssd1 vssd1 vccd1 vccd1 hold504/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3503_ _3504_/CLK _3503_/D _2997_/Y vssd1 vssd1 vccd1 vccd1 _3503_/Q sky130_fd_sc_hd__dfrtp_1
X_3434_ _3434_/CLK _3434_/D vssd1 vssd1 vccd1 vccd1 _3434_/Q sky130_fd_sc_hd__dfxtp_1
Xhold537 _2815_/X vssd1 vssd1 vccd1 vccd1 _3338_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 _3335_/Q vssd1 vssd1 vccd1 vccd1 hold548/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 _2837_/X vssd1 vssd1 vccd1 vccd1 _3368_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1695_ _1697_/B _1697_/C _1697_/A vssd1 vssd1 vccd1 vccd1 _1695_/X sky130_fd_sc_hd__or3b_1
XANTENNA__2026__S1 _2195_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _3424_/CLK _3365_/D vssd1 vssd1 vccd1 vccd1 _3365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _3484_/CLK _3296_/D vssd1 vssd1 vccd1 vccd1 _3296_/Q sky130_fd_sc_hd__dfxtp_1
X_2316_ _2316_/A _2316_/B vssd1 vssd1 vccd1 vccd1 _2316_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2247_ _2249_/A _3464_/Q _3463_/Q _2246_/X hold846/X vssd1 vssd1 vccd1 vccd1 _2247_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_79_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2178_ _3591_/Q _2578_/B vssd1 vssd1 vccd1 vccd1 _2178_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2721__S _2728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1917__A1 _2546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2017__S1 _2219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput57 _3654_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_12
Xoutput46 _2571_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_12
XANTENNA_fanout96_A _3483_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2631__S _2633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2581__A1 _2801_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3150_ _3550_/CLK _3150_/D _2914_/Y vssd1 vssd1 vccd1 vccd1 _3150_/Q sky130_fd_sc_hd__dfrtp_1
X_3081_ _3090_/A vssd1 vssd1 vccd1 vccd1 _3081_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_27_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2101_ _2061_/X _2090_/A _2100_/X vssd1 vssd1 vccd1 vccd1 _2101_/Y sky130_fd_sc_hd__a21oi_2
X_2032_ _2144_/C _2316_/A _2023_/Y vssd1 vssd1 vccd1 vccd1 _2032_/Y sky130_fd_sc_hd__o21ai_1
X_2934_ _3122_/A vssd1 vssd1 vccd1 vccd1 _2934_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2495__S1 _1912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2865_ hold516/X _2105_/A _2870_/S vssd1 vssd1 vccd1 vccd1 _2865_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1946__A _2546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1816_ _1886_/A _1816_/B vssd1 vssd1 vccd1 vccd1 _1816_/Y sky130_fd_sc_hd__nor2_1
X_2796_ hold280/X _2806_/A1 _2799_/S vssd1 vssd1 vccd1 vccd1 _2796_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold301 _3311_/Q vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 _3264_/Q vssd1 vssd1 vccd1 vccd1 hold334/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 _3594_/Q vssd1 vssd1 vccd1 vccd1 hold323/X sky130_fd_sc_hd__dlygate4sd3_1
X_1747_ _1811_/S _1747_/B _1769_/B vssd1 vssd1 vccd1 vccd1 _1747_/X sky130_fd_sc_hd__or3_1
Xhold312 _3330_/Q vssd1 vssd1 vccd1 vccd1 hold312/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold345 _3246_/Q vssd1 vssd1 vccd1 vccd1 hold345/X sky130_fd_sc_hd__dlygate4sd3_1
X_1678_ _3601_/Q hold59/X hold65/X vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__mux2_1
Xhold367 _2757_/X vssd1 vssd1 vccd1 vccd1 _3286_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 _2660_/X vssd1 vssd1 vccd1 vccd1 _3201_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 _3219_/Q vssd1 vssd1 vccd1 vccd1 hold378/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3417_ _3516_/CLK _3417_/D vssd1 vssd1 vccd1 vccd1 _3417_/Q sky130_fd_sc_hd__dfxtp_1
Xhold389 _2703_/X vssd1 vssd1 vccd1 vccd1 _3239_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3348_ _3550_/CLK _3348_/D _2923_/Y vssd1 vssd1 vccd1 vccd1 _3348_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 _2239_/X vssd1 vssd1 vccd1 vccd1 _2240_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 _3521_/Q vssd1 vssd1 vccd1 vccd1 _1891_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 _2363_/A vssd1 vssd1 vccd1 vccd1 _2385_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ _3484_/CLK _3279_/D vssd1 vssd1 vccd1 vccd1 _3279_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1034 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 hold125/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1045 _3549_/Q vssd1 vssd1 vccd1 vccd1 hold948/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2716__S _2718_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2451__S _2546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold890 _2193_/Y vssd1 vssd1 vccd1 vccd1 hold890/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2626__S _2633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2650_ _2104_/B hold686/X _2654_/S vssd1 vssd1 vccd1 vccd1 _2650_/X sky130_fd_sc_hd__mux2_1
X_1601_ _1808_/D vssd1 vssd1 vccd1 vccd1 _1601_/Y sky130_fd_sc_hd__inv_2
X_2581_ hold423/X _2801_/A1 _2589_/S vssd1 vssd1 vccd1 vccd1 _2581_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3202_ _3333_/CLK _3202_/D vssd1 vssd1 vccd1 vccd1 _3202_/Q sky130_fd_sc_hd__dfxtp_1
X_3133_ _3326_/CLK _3133_/D vssd1 vssd1 vccd1 vccd1 _3133_/Q sky130_fd_sc_hd__dfxtp_1
X_3064_ _3067_/A vssd1 vssd1 vccd1 vccd1 _3064_/Y sky130_fd_sc_hd__inv_2
X_2015_ hold237/X hold241/X hold210/X hold243/X _2045_/S0 _2045_/S1 vssd1 vssd1 vccd1
+ vccd1 _2015_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2917_ _3049_/A vssd1 vssd1 vccd1 vccd1 _2917_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2793__A1 _2803_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2848_ _2355_/B hold658/X _2849_/S vssd1 vssd1 vccd1 vccd1 _2848_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2779_ hold40/X hold30/X _2779_/S vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__mux2_1
XFILLER_0_5_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold120 input28/X vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold131 _3245_/Q vssd1 vssd1 vccd1 vccd1 hold131/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold153 _1661_/X vssd1 vssd1 vccd1 vccd1 _1665_/S sky130_fd_sc_hd__clkbuf_2
Xhold142 _3290_/Q vssd1 vssd1 vccd1 vccd1 hold142/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 _3131_/Q vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _2802_/X vssd1 vssd1 vccd1 vccd1 _3326_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _2680_/X vssd1 vssd1 vccd1 vccd1 _3218_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 _2727_/X vssd1 vssd1 vccd1 vccd1 _3260_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2775__A1 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2702_ _2804_/A1 hold194/X _2707_/S vssd1 vssd1 vccd1 vccd1 _2702_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2633_ _2356_/B hold634/X _2633_/S vssd1 vssd1 vccd1 vccd1 _2633_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2104__B _2104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2564_ _2574_/A _2564_/B vssd1 vssd1 vccd1 vccd1 _2564_/X sky130_fd_sc_hd__and2_2
XANTENNA__2527__A1 _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2495_ _3176_/Q _3425_/Q _3416_/Q _3158_/Q _1918_/B _1912_/B vssd1 vssd1 vccd1 vccd1
+ _2495_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_4_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3116_ _3129_/A vssd1 vssd1 vccd1 vccd1 _3116_/Y sky130_fd_sc_hd__inv_2
X_3047_ _3049_/A vssd1 vssd1 vccd1 vccd1 _3047_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_73_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2757__A1 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout92 hold909/X vssd1 vssd1 vccd1 vccd1 _2222_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout70 _2106_/X vssd1 vssd1 vccd1 vccd1 _2360_/B sky130_fd_sc_hd__buf_4
Xfanout81 hold311/X vssd1 vssd1 vccd1 vccd1 _2121_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1747__C _1769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2280_ _2271_/B _2281_/B _2279_/Y vssd1 vssd1 vccd1 vccd1 _2280_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_19_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1995_ _3249_/Q _3321_/Q _3312_/Q _3303_/Q _2049_/S0 _2219_/A vssd1 vssd1 vccd1 vccd1
+ _1995_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_7_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2616_ _2098_/S hold772/X _2623_/S vssd1 vssd1 vccd1 vccd1 _2616_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout109_A hold120/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3596_ _3600_/CLK _3596_/D _3087_/Y vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dfrtp_1
X_2547_ _2543_/X _2546_/X _3518_/Q vssd1 vssd1 vccd1 vccd1 _2547_/X sky130_fd_sc_hd__mux2_1
X_2478_ _3637_/Q _2510_/A _2475_/X _2477_/X _2510_/B vssd1 vssd1 vccd1 vccd1 _2478_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2684__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2531__S0 _1918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2724__S _2728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2739__A1 _2406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1650__A1 hold75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1780_ _2092_/A _3552_/Q vssd1 vssd1 vccd1 vccd1 _1784_/B sky130_fd_sc_hd__or2_1
XFILLER_0_37_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold708 _3181_/Q vssd1 vssd1 vccd1 vccd1 hold708/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold719 _2866_/X vssd1 vssd1 vccd1 vccd1 _3398_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3450_ _3632_/CLK hold6/X _2944_/Y vssd1 vssd1 vccd1 vccd1 _3450_/Q sky130_fd_sc_hd__dfrtp_1
X_2401_ _2401_/A hold98/X hold95/X vssd1 vssd1 vccd1 vccd1 _3583_/D sky130_fd_sc_hd__and3_1
X_3381_ _3600_/CLK _3381_/D _2929_/Y vssd1 vssd1 vccd1 vccd1 _3381_/Q sky130_fd_sc_hd__dfrtp_1
X_2332_ _3383_/Q _2267_/X hold854/X vssd1 vssd1 vccd1 vccd1 _2332_/X sky130_fd_sc_hd__o21ba_1
X_2263_ _1558_/Y hold806/X _1593_/Y hold80/X vssd1 vssd1 vccd1 vccd1 _2263_/X sky130_fd_sc_hd__a22o_1
X_2194_ _2219_/A _2221_/B _2211_/A vssd1 vssd1 vccd1 vccd1 _2194_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__2666__A0 _2406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1641__A1 _2399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1978_ hold780/X _1977_/Y _2000_/S vssd1 vssd1 vccd1 vccd1 _1978_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3648_ _3655_/A vssd1 vssd1 vccd1 vccd1 _3648_/X sky130_fd_sc_hd__buf_1
X_3579_ _3579_/CLK _3579_/D vssd1 vssd1 vccd1 vccd1 _3579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3333_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__clkbuf_2
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2629__S _2633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2648__A0 _2109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2950_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2950_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2881_ _2891_/B _2881_/B vssd1 vssd1 vccd1 vccd1 _2890_/S sky130_fd_sc_hd__nand2_8
X_1901_ _2891_/A vssd1 vssd1 vccd1 vccd1 _1901_/Y sky130_fd_sc_hd__inv_2
X_1832_ _3543_/Q hold844/X _1835_/S vssd1 vssd1 vccd1 vccd1 _1832_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_40_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1763_ _1811_/S _3557_/Q _1769_/B vssd1 vssd1 vccd1 vccd1 _1763_/X sky130_fd_sc_hd__or3_1
Xhold527 _2899_/X vssd1 vssd1 vccd1 vccd1 _3428_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 _3397_/Q vssd1 vssd1 vccd1 vccd1 hold516/X sky130_fd_sc_hd__dlygate4sd3_1
X_1694_ hold908/X _1697_/C _1697_/A vssd1 vssd1 vccd1 vccd1 _1694_/X sky130_fd_sc_hd__o21a_1
Xhold505 _2652_/X vssd1 vssd1 vccd1 vccd1 _3196_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3502_ _3610_/CLK _3502_/D _2996_/Y vssd1 vssd1 vccd1 vccd1 _3502_/Q sky130_fd_sc_hd__dfrtp_1
Xhold538 _3421_/Q vssd1 vssd1 vccd1 vccd1 hold538/X sky130_fd_sc_hd__dlygate4sd3_1
X_3433_ _3433_/CLK _3433_/D vssd1 vssd1 vccd1 vccd1 _3433_/Q sky130_fd_sc_hd__dfxtp_1
Xhold549 _2812_/X vssd1 vssd1 vccd1 vccd1 _3335_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _3413_/CLK _3364_/D vssd1 vssd1 vccd1 vccd1 _3364_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _3484_/CLK _3295_/D vssd1 vssd1 vccd1 vccd1 _3295_/Q sky130_fd_sc_hd__dfxtp_1
X_2315_ _2315_/A1 _2018_/X _2019_/X _2014_/X _1774_/X vssd1 vssd1 vccd1 vccd1 _2316_/B
+ sky130_fd_sc_hd__o221ai_2
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2639__A0 _2104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2246_ _2248_/A _3469_/Q _3468_/Q _3467_/Q vssd1 vssd1 vccd1 vccd1 _2246_/X sky130_fd_sc_hd__and4_1
XFILLER_0_79_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2177_ _2177_/A _2177_/B _2800_/A vssd1 vssd1 vccd1 vccd1 _3488_/D sky130_fd_sc_hd__and3_1
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput47 _2573_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_12
Xoutput58 _2470_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_12
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2878__A0 _2357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2973__A _3124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1755__C _1769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2030__A1 _2036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2333__A2 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3080_ _3090_/A vssd1 vssd1 vccd1 vccd1 _3080_/Y sky130_fd_sc_hd__inv_2
X_2100_ _2064_/B _2078_/X _2085_/X _2064_/A _2067_/B vssd1 vssd1 vccd1 vccd1 _2100_/X
+ sky130_fd_sc_hd__a221o_1
X_2031_ _2315_/A1 _2029_/X _2030_/Y _2025_/Y vssd1 vssd1 vccd1 vccd1 _2316_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_43_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2933_ _3129_/A vssd1 vssd1 vccd1 vccd1 _2933_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2822__S _2829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2864_ hold514/X _2109_/B _2870_/S vssd1 vssd1 vccd1 vccd1 _2864_/X sky130_fd_sc_hd__mux2_1
X_2795_ hold332/X _2805_/A1 _2799_/S vssd1 vssd1 vccd1 vccd1 _2795_/X sky130_fd_sc_hd__mux2_1
X_1815_ _1886_/B _1810_/Y _1814_/B vssd1 vssd1 vccd1 vccd1 _1815_/X sky130_fd_sc_hd__a21o_1
X_1746_ hold921/X _2387_/C _1745_/X vssd1 vssd1 vccd1 vccd1 _1746_/X sky130_fd_sc_hd__o21a_1
Xhold302 _2785_/X vssd1 vssd1 vccd1 vccd1 _3311_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 _2733_/X vssd1 vssd1 vccd1 vccd1 _3264_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 _2806_/X vssd1 vssd1 vccd1 vccd1 _3330_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 _3228_/Q vssd1 vssd1 vccd1 vccd1 hold324/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 _3252_/Q vssd1 vssd1 vccd1 vccd1 hold357/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 _2712_/X vssd1 vssd1 vccd1 vccd1 _3246_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 _3313_/Q vssd1 vssd1 vccd1 vccd1 hold368/X sky130_fd_sc_hd__dlygate4sd3_1
X_1677_ _2289_/A hold64/X vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__nor2_1
X_3416_ _3431_/CLK _3416_/D vssd1 vssd1 vccd1 vccd1 _3416_/Q sky130_fd_sc_hd__dfxtp_1
Xhold379 _2681_/X vssd1 vssd1 vccd1 vccd1 _3219_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3347_ _3635_/CLK _3347_/D _2922_/Y vssd1 vssd1 vccd1 vccd1 _3347_/Q sky130_fd_sc_hd__dfstp_1
Xhold1002 _3531_/Q vssd1 vssd1 vccd1 vccd1 _1847_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold1024 _3578_/Q vssd1 vssd1 vccd1 vccd1 hold465/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1013 _1898_/X vssd1 vssd1 vccd1 vccd1 _3521_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3278_ _3484_/CLK _3278_/D vssd1 vssd1 vccd1 vccd1 _3278_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1046 _3497_/Q vssd1 vssd1 vccd1 vccd1 hold997/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__dlygate4sd3_1
X_2229_ _2259_/A _2259_/B _2240_/A vssd1 vssd1 vccd1 vccd1 _2230_/B sky130_fd_sc_hd__and3_1
XFILLER_0_82_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2260__A1 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold880 _3460_/Q vssd1 vssd1 vccd1 vccd1 _2272_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 _2196_/Y vssd1 vssd1 vccd1 vccd1 _3483_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1600_ _1825_/A vssd1 vssd1 vccd1 vccd1 _1600_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_22_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2580_ _2790_/A _2719_/A vssd1 vssd1 vccd1 vccd1 _2589_/S sky130_fd_sc_hd__nor2_4
XFILLER_0_10_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3201_ _3332_/CLK _3201_/D vssd1 vssd1 vccd1 vccd1 _3201_/Q sky130_fd_sc_hd__dfxtp_1
X_3132_ _3320_/CLK _3132_/D vssd1 vssd1 vccd1 vccd1 _3132_/Q sky130_fd_sc_hd__dfxtp_1
X_3063_ _3069_/A vssd1 vssd1 vccd1 vccd1 _3063_/Y sky130_fd_sc_hd__inv_2
X_2014_ _2036_/S _2014_/B vssd1 vssd1 vccd1 vccd1 _2014_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2916_ _3054_/A vssd1 vssd1 vccd1 vccd1 _2916_/Y sky130_fd_sc_hd__inv_2
X_2847_ _2357_/B hold546/X _2849_/S vssd1 vssd1 vccd1 vccd1 _2847_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2778_ hold239/X _2808_/A1 _2779_/S vssd1 vssd1 vccd1 vccd1 _2778_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold110 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 input12/A sky130_fd_sc_hd__dlygate4sd3_1
X_1729_ _1581_/Y _3452_/Q _1711_/Y _1719_/Y _1723_/Y vssd1 vssd1 vccd1 vccd1 _1739_/C
+ sky130_fd_sc_hd__o2111ai_2
Xhold121 _1670_/X vssd1 vssd1 vccd1 vccd1 _3605_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 _2711_/X vssd1 vssd1 vccd1 vccd1 _3245_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 _2762_/X vssd1 vssd1 vccd1 vccd1 _3290_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 _3236_/Q vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _1662_/X vssd1 vssd1 vccd1 vccd1 _3610_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _3283_/Q vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 _2582_/X vssd1 vssd1 vccd1 vccd1 _3131_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 _3637_/Q vssd1 vssd1 vccd1 vccd1 _1768_/S sky130_fd_sc_hd__buf_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1631__S hold12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2727__S _2728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2701_ _2803_/A1 hold316/X _2707_/S vssd1 vssd1 vccd1 vccd1 _2701_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2632_ _2355_/B hold648/X _2633_/S vssd1 vssd1 vccd1 vccd1 _2632_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2563_ _3451_/Q _2510_/B _2559_/X _2562_/X vssd1 vssd1 vccd1 vccd1 _2564_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2401__A _2401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2494_ _3407_/Q _3398_/Q _3389_/Q _3434_/Q _2532_/S0 _2532_/S1 vssd1 vssd1 vccd1
+ vccd1 _2494_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2547__S _3518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3115_ _3127_/A vssd1 vssd1 vccd1 vccd1 _3115_/Y sky130_fd_sc_hd__inv_2
X_3046_ _3049_/A vssd1 vssd1 vccd1 vccd1 _3046_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout71_A _2101_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2014__A_N _2036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1597__A _2144_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout82 hold477/X vssd1 vssd1 vccd1 vccd1 _2546_/S sky130_fd_sc_hd__buf_6
Xfanout71 _2101_/Y vssd1 vssd1 vccd1 vccd1 _2105_/A sky130_fd_sc_hd__buf_4
Xfanout93 _2195_/A1 vssd1 vssd1 vccd1 vccd1 _2045_/S1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1763__C _1769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3576_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2693__A1 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1994_ _3294_/Q _3285_/Q _3276_/Q _3267_/Q _2049_/S0 _2195_/A1 vssd1 vssd1 vccd1
+ vccd1 _1994_/X sky130_fd_sc_hd__mux4_1
XANTENNA__1657__D input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2115__B _2383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2615_ _2358_/B hold650/X _2623_/S vssd1 vssd1 vccd1 vccd1 _2615_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3595_ _3607_/CLK _3595_/D _3086_/Y vssd1 vssd1 vccd1 vccd1 _3595_/Q sky130_fd_sc_hd__dfrtp_1
X_2546_ _2545_/X _2544_/X _2546_/S vssd1 vssd1 vccd1 vccd1 _2546_/X sky130_fd_sc_hd__mux2_1
X_2477_ _3623_/Q hold11/A hold52/A _3614_/Q _2476_/X vssd1 vssd1 vccd1 vccd1 _2477_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3029_ _3032_/A vssd1 vssd1 vccd1 vccd1 _3029_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2531__S1 _1912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2047__S0 _3483_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2976__A _3124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2675__A1 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2650__S _2654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold709 _2635_/X vssd1 vssd1 vccd1 vccd1 _3181_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2038__S0 _2221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2400_ _2400_/A hold98/X hold95/X vssd1 vssd1 vccd1 vccd1 _3582_/D sky130_fd_sc_hd__and3_1
X_3380_ _3600_/CLK _3380_/D _2928_/Y vssd1 vssd1 vccd1 vccd1 _3380_/Q sky130_fd_sc_hd__dfrtp_1
X_2331_ _1923_/A hold860/X _3581_/Q vssd1 vssd1 vccd1 vccd1 _2331_/X sky130_fd_sc_hd__o21ba_1
X_2262_ hold67/X _2270_/A vssd1 vssd1 vccd1 vccd1 _2267_/D sky130_fd_sc_hd__xnor2_1
X_2193_ _2193_/A _2193_/B vssd1 vssd1 vccd1 vccd1 _2193_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2825__S _2829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_47_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout121_A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1977_ _1977_/A vssd1 vssd1 vccd1 vccd1 _1977_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3647_ _3655_/A vssd1 vssd1 vccd1 vccd1 _3647_/X sky130_fd_sc_hd__buf_1
XFILLER_0_11_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3578_ _3579_/CLK input1/X vssd1 vssd1 vccd1 vccd1 _3578_/Q sky130_fd_sc_hd__dfxtp_1
X_2529_ _3188_/Q _3341_/Q _3170_/Q _3146_/Q _2532_/S0 _1943_/A vssd1 vssd1 vccd1 vccd1
+ _2529_/X sky130_fd_sc_hd__mux4_1
Xhold14 wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__clkbuf_4
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2593__A0 _2358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2896__A1 _2104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1769__B _1769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2880_ _2356_/B hold690/X _2880_/S vssd1 vssd1 vccd1 vccd1 _2880_/X sky130_fd_sc_hd__mux2_1
X_1900_ _1902_/A _1905_/B vssd1 vssd1 vccd1 vccd1 _2891_/A sky130_fd_sc_hd__nor2_2
X_1831_ hold838/X _3543_/Q _1835_/S vssd1 vssd1 vccd1 vccd1 _1831_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1762_ hold969/X _2387_/C _1761_/X vssd1 vssd1 vccd1 vccd1 _1762_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_4_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold517 _2865_/X vssd1 vssd1 vccd1 vccd1 _3397_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold506 _3399_/Q vssd1 vssd1 vccd1 vccd1 hold506/X sky130_fd_sc_hd__dlygate4sd3_1
X_1693_ _1698_/A _1698_/B vssd1 vssd1 vccd1 vccd1 _1697_/C sky130_fd_sc_hd__or2_2
X_3501_ _3638_/CLK _3501_/D _2995_/Y vssd1 vssd1 vccd1 vccd1 _3501_/Q sky130_fd_sc_hd__dfrtp_1
Xhold539 _2892_/X vssd1 vssd1 vccd1 vccd1 _3421_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3432_ _3432_/CLK _3432_/D vssd1 vssd1 vccd1 vccd1 _3432_/Q sky130_fd_sc_hd__dfxtp_1
Xhold528 _3353_/Q vssd1 vssd1 vccd1 vccd1 hold528/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3424_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3363_ _3413_/CLK _3363_/D vssd1 vssd1 vccd1 vccd1 _3363_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2431__S0 _1918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _3321_/CLK _3294_/D vssd1 vssd1 vccd1 vccd1 _3294_/Q sky130_fd_sc_hd__dfxtp_1
X_2314_ _2314_/A _2314_/B vssd1 vssd1 vccd1 vccd1 _2323_/A sky130_fd_sc_hd__nand2_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2245_ _3472_/Q _2205_/B _2244_/X _2183_/Y _2211_/A vssd1 vssd1 vccd1 vccd1 _2245_/X
+ sky130_fd_sc_hd__a221o_1
X_2176_ _2176_/A _2578_/B vssd1 vssd1 vccd1 vccd1 _2800_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_79_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2811__A1 _2358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput48 _3646_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_12
Xoutput59 _3655_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_12
XANTENNA__1634__S hold12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2465__S _2546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2802__A1 _2802_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2522__B1_N hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2869__A1 _2355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2030_ _2036_/S _2026_/X _2315_/A1 vssd1 vssd1 vccd1 vccd1 _2030_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_43_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2932_ _3090_/A vssd1 vssd1 vccd1 vccd1 _2932_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2863_ hold614/X _2098_/S _2870_/S vssd1 vssd1 vccd1 vccd1 _2863_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2404__A hold87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1814_ _1886_/B _1814_/B vssd1 vssd1 vccd1 vccd1 _1814_/Y sky130_fd_sc_hd__nor2_1
X_2794_ hold169/X _2804_/A1 _2799_/S vssd1 vssd1 vccd1 vccd1 _2794_/X sky130_fd_sc_hd__mux2_1
X_1745_ _1811_/S _3566_/Q _1769_/B vssd1 vssd1 vccd1 vccd1 _1745_/X sky130_fd_sc_hd__or3_1
XFILLER_0_13_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2021__A2 _2144_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold303 _3213_/Q vssd1 vssd1 vccd1 vccd1 hold303/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 _2691_/X vssd1 vssd1 vccd1 vccd1 _3228_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 _3284_/Q vssd1 vssd1 vccd1 vccd1 hold314/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 _3300_/Q vssd1 vssd1 vccd1 vccd1 hold336/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 _2718_/X vssd1 vssd1 vccd1 vccd1 _3252_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 _3273_/Q vssd1 vssd1 vccd1 vccd1 hold347/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 _2787_/X vssd1 vssd1 vccd1 vccd1 _3313_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1676_ _2421_/B hold63/X vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__nand2_1
X_3415_ _3424_/CLK _3415_/D vssd1 vssd1 vccd1 vccd1 _3415_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3346_ _3635_/CLK _3346_/D _2921_/Y vssd1 vssd1 vccd1 vccd1 _3346_/Q sky130_fd_sc_hd__dfrtp_2
Xhold1003 _1870_/X vssd1 vssd1 vccd1 vccd1 _3531_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1014 _3522_/Q vssd1 vssd1 vccd1 vccd1 _1892_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1025 _3297_/Q vssd1 vssd1 vccd1 vccd1 _2769_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_3277_ _3322_/CLK _3277_/D vssd1 vssd1 vccd1 vccd1 _3277_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1036 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 input4/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1047 _3511_/Q vssd1 vssd1 vccd1 vccd1 hold822/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2228_ _2363_/A _2228_/B _2228_/C vssd1 vssd1 vccd1 vccd1 _2240_/A sky130_fd_sc_hd__and3b_1
X_2159_ _3522_/Q _2159_/B vssd1 vssd1 vccd1 vccd1 _2161_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1629__S hold12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold881 _2276_/X vssd1 vssd1 vccd1 vccd1 _3460_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold870 _2238_/Y vssd1 vssd1 vccd1 vccd1 _3474_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 _3572_/Q vssd1 vssd1 vccd1 vccd1 _1700_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2720__A0 _2801_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2787__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3055__A _3057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3200_ _3326_/CLK _3200_/D vssd1 vssd1 vccd1 vccd1 _3200_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2711__A0 _2802_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3131_ _3408_/CLK _3131_/D vssd1 vssd1 vccd1 vccd1 _3131_/Q sky130_fd_sc_hd__dfxtp_1
X_3062_ _3069_/A vssd1 vssd1 vccd1 vccd1 _3062_/Y sky130_fd_sc_hd__inv_2
X_2013_ hold190/X hold214/X hold194/X hold206/X _2045_/S0 _2045_/S1 vssd1 vssd1 vccd1
+ vccd1 _2014_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_77_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2915_ _3054_/A vssd1 vssd1 vccd1 vccd1 _2915_/Y sky130_fd_sc_hd__inv_2
X_2846_ _2106_/X hold776/X _2849_/S vssd1 vssd1 vccd1 vccd1 _2846_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold100 _3638_/Q vssd1 vssd1 vccd1 vccd1 _1767_/S sky130_fd_sc_hd__buf_2
X_2777_ hold384/X _2807_/A1 _2779_/S vssd1 vssd1 vccd1 vccd1 _2777_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_73 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1728_ _1885_/S hold338/X _1713_/Y _1715_/Y _1728_/D1 vssd1 vssd1 vccd1 vccd1 _1739_/B
+ sky130_fd_sc_hd__o2111ai_2
Xhold144 _3614_/Q vssd1 vssd1 vccd1 vccd1 _1568_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 _1623_/C vssd1 vssd1 vccd1 vccd1 _1655_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 input20/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 _3263_/Q vssd1 vssd1 vccd1 vccd1 hold133/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 _2700_/X vssd1 vssd1 vccd1 vccd1 _3236_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1659_ hold62/X _1659_/B _1659_/C vssd1 vssd1 vccd1 vccd1 _2421_/A sky130_fd_sc_hd__and3b_2
Xhold155 _3292_/Q vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 _2754_/X vssd1 vssd1 vccd1 vccd1 _3283_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _3278_/Q vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _1619_/X vssd1 vssd1 vccd1 vccd1 _3637_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2702__A0 _2804_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _3329_/CLK _3329_/D vssd1 vssd1 vccd1 vccd1 _3329_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2743__S _2749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2769__A0 hold30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2219__A _2219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2653__S _2654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2700_ _2802_/A1 hold176/X _2707_/S vssd1 vssd1 vccd1 vccd1 _2700_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_27_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2631_ _2357_/B hold630/X _2633_/S vssd1 vssd1 vccd1 vccd1 _2631_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2562_ hold80/A hold11/A vssd1 vssd1 vccd1 vccd1 _2562_/X sky130_fd_sc_hd__or2_1
XFILLER_0_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2493_ _3185_/Q _3338_/Q _3167_/Q _3143_/Q _1944_/B _1943_/A vssd1 vssd1 vccd1 vccd1
+ _2493_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2828__S _2829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3114_ _3129_/A vssd1 vssd1 vccd1 vccd1 _3114_/Y sky130_fd_sc_hd__inv_2
X_3045_ _3054_/A vssd1 vssd1 vccd1 vccd1 _3045_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1671__A0 _2399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2829_ hold508/X _2356_/B _2829_/S vssd1 vssd1 vccd1 vccd1 _2829_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1642__S hold12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout72 _2097_/X vssd1 vssd1 vccd1 vccd1 _2358_/B sky130_fd_sc_hd__buf_4
Xfanout83 _2532_/S1 vssd1 vssd1 vccd1 vccd1 _1943_/A sky130_fd_sc_hd__clkbuf_8
Xfanout94 _2195_/A1 vssd1 vssd1 vccd1 vccd1 _2219_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2221__B _2221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2648__S _2654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_47_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1993_ _1991_/X _1992_/X _2036_/S vssd1 vssd1 vccd1 vccd1 _1993_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2614_ _2810_/B _2881_/B vssd1 vssd1 vccd1 vccd1 _2623_/S sky130_fd_sc_hd__nand2_4
X_3594_ _3594_/CLK _3594_/D _3085_/Y vssd1 vssd1 vccd1 vccd1 _3594_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2905__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2545_ _3189_/Q _3342_/Q _3171_/Q _3147_/Q _1944_/B _1943_/A vssd1 vssd1 vccd1 vccd1
+ _2545_/X sky130_fd_sc_hd__mux4_1
X_2476_ _3514_/Q _2507_/C _2572_/A vssd1 vssd1 vccd1 vccd1 _2476_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3028_ _3032_/A vssd1 vssd1 vccd1 vccd1 _3028_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_65_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1947__A1 _3518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold111_A _1623_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1637__S hold12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2047__S1 _2195_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2468__S _2546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2038__S1 _2219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2330_ _2144_/D _2327_/X hold876/X vssd1 vssd1 vccd1 vccd1 _2330_/X sky130_fd_sc_hd__a21o_1
X_2261_ _3632_/Q _3460_/Q vssd1 vssd1 vccd1 vccd1 _2261_/Y sky130_fd_sc_hd__xnor2_1
X_2192_ _2186_/X _2243_/B _2222_/A _2193_/B vssd1 vssd1 vccd1 vccd1 _3485_/D sky130_fd_sc_hd__a2bb2o_1
XANTENNA__2407__A hold59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2841__S _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1976_ _2225_/A _1971_/X _1975_/X vssd1 vssd1 vccd1 vccd1 _1977_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3646_ _3655_/A vssd1 vssd1 vccd1 vccd1 _3646_/X sky130_fd_sc_hd__buf_1
XANTENNA_fanout114_A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3577_ _3627_/CLK _3577_/D _3070_/Y vssd1 vssd1 vccd1 vccd1 _3577_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2528_ _3410_/Q _3401_/Q _3392_/Q _3437_/Q _1944_/B _2532_/S1 vssd1 vssd1 vccd1 vccd1
+ _2528_/X sky130_fd_sc_hd__mux4_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__buf_1
X_2459_ _3513_/Q _2507_/C _2572_/A vssd1 vssd1 vccd1 vccd1 _2459_/X sky130_fd_sc_hd__o21a_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__buf_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1960__S0 _2045_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1769__C _2383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1830_ hold811/X _3544_/Q _1835_/S vssd1 vssd1 vccd1 vccd1 _1830_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_37_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1761_ _3148_/Q _1761_/B _1769_/B vssd1 vssd1 vccd1 vccd1 _1761_/X sky130_fd_sc_hd__or3_1
XFILLER_0_4_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2584__A1 _2804_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3500_ _3576_/CLK _3500_/D _2994_/Y vssd1 vssd1 vccd1 vccd1 _3500_/Q sky130_fd_sc_hd__dfrtp_1
Xhold518 _3423_/Q vssd1 vssd1 vccd1 vccd1 hold518/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold507 _2867_/X vssd1 vssd1 vccd1 vccd1 _3399_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1692_ _1700_/A _1700_/B vssd1 vssd1 vccd1 vccd1 _1698_/B sky130_fd_sc_hd__or2_1
X_3431_ _3431_/CLK _3431_/D vssd1 vssd1 vccd1 vccd1 _3431_/Q sky130_fd_sc_hd__dfxtp_1
Xhold529 _2821_/X vssd1 vssd1 vccd1 vccd1 _3353_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ _3431_/CLK _3362_/D vssd1 vssd1 vccd1 vccd1 _3362_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2431__S1 _1912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2313_ _1564_/Y _1977_/A _1988_/A _2312_/X vssd1 vssd1 vccd1 vccd1 _2314_/B sky130_fd_sc_hd__o31a_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _3322_/CLK _3293_/D vssd1 vssd1 vccd1 vccd1 _3293_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ _2708_/A _2241_/B _2242_/X _2243_/X vssd1 vssd1 vccd1 vccd1 _2244_/X sky130_fd_sc_hd__o211a_1
X_2175_ _2176_/A _2578_/B vssd1 vssd1 vccd1 vccd1 _2177_/B sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3322_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1959_ hold403/X hold409/X hold437/X hold445/X _2045_/S0 _2045_/S1 vssd1 vssd1 vccd1
+ vccd1 _1959_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_43_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3629_ _3633_/CLK _3629_/D _3120_/Y vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__dfstp_1
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput38 _2395_/X vssd1 vssd1 vccd1 vccd1 uart_irq sky130_fd_sc_hd__buf_12
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput49 _3647_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_12
XANTENNA__2746__S _2749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2931_ _3122_/A vssd1 vssd1 vccd1 vccd1 _2931_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_84_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2862_ hold502/X _2358_/B _2870_/S vssd1 vssd1 vccd1 vccd1 _2862_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2793_ hold372/X _2803_/A1 _2799_/S vssd1 vssd1 vccd1 vccd1 _2793_/X sky130_fd_sc_hd__mux2_1
X_1813_ _2383_/A _1813_/B vssd1 vssd1 vccd1 vccd1 _1814_/B sky130_fd_sc_hd__or2_1
XFILLER_0_25_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1744_ _1886_/A _2383_/A _1886_/B vssd1 vssd1 vccd1 vccd1 _1769_/B sky130_fd_sc_hd__or3_4
Xhold326 _3442_/Q vssd1 vssd1 vccd1 vccd1 _1726_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold304 _2673_/X vssd1 vssd1 vccd1 vccd1 _3213_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 _2755_/X vssd1 vssd1 vccd1 vccd1 _3284_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 _2773_/X vssd1 vssd1 vccd1 vccd1 _3300_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 _2743_/X vssd1 vssd1 vccd1 vccd1 _3273_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold359 _3250_/Q vssd1 vssd1 vccd1 vccd1 hold359/X sky130_fd_sc_hd__dlygate4sd3_1
X_3414_ _3579_/CLK _3414_/D vssd1 vssd1 vccd1 vccd1 _3414_/Q sky130_fd_sc_hd__dfxtp_1
X_1675_ _2421_/B hold63/A vssd1 vssd1 vccd1 vccd1 _1675_/X sky130_fd_sc_hd__and2_1
XFILLER_0_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3345_ _3594_/CLK _3345_/D _2920_/Y vssd1 vssd1 vccd1 vccd1 _3345_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1004 hold1055/X vssd1 vssd1 vccd1 vccd1 _1850_/A sky130_fd_sc_hd__buf_1
X_3276_ _3321_/CLK _3276_/D vssd1 vssd1 vccd1 vccd1 _3276_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1015 _1894_/X vssd1 vssd1 vccd1 vccd1 _3522_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1026 _3315_/Q vssd1 vssd1 vccd1 vccd1 _2789_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 hold116/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1037 _1610_/X vssd1 vssd1 vccd1 vccd1 _1611_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ _2227_/A _2227_/B vssd1 vssd1 vccd1 vccd1 _2227_/X sky130_fd_sc_hd__and2_1
XFILLER_0_84_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2158_ _2157_/Y _2157_/A _2158_/S vssd1 vssd1 vccd1 vccd1 _3492_/D sky130_fd_sc_hd__mux2_1
X_2089_ _2059_/Y _2068_/Y _2077_/Y _2084_/Y _2092_/A _2058_/C vssd1 vssd1 vccd1 vccd1
+ _2090_/B sky130_fd_sc_hd__mux4_2
XFILLER_0_48_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2796__A1 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1923__C_N _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout94_A _2195_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold871 _3576_/Q vssd1 vssd1 vccd1 vccd1 hold871/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold882 _3583_/Q vssd1 vssd1 vccd1 vccd1 hold882/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold860 _3384_/Q vssd1 vssd1 vccd1 vccd1 hold860/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 _1700_/Y vssd1 vssd1 vccd1 vccd1 hold893/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3130_ _3329_/CLK _3130_/D vssd1 vssd1 vccd1 vccd1 _3130_/Q sky130_fd_sc_hd__dfxtp_1
X_3061_ _3061_/A vssd1 vssd1 vccd1 vccd1 _3061_/Y sky130_fd_sc_hd__inv_2
X_2012_ hold796/X _2011_/Y _2055_/S vssd1 vssd1 vccd1 vccd1 _2012_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2778__A1 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2914_ _3129_/A vssd1 vssd1 vccd1 vccd1 _2914_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2845_ _2104_/B hold728/X _2849_/S vssd1 vssd1 vccd1 vccd1 _2845_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2776_ hold286/X _2806_/A1 _2779_/S vssd1 vssd1 vccd1 vccd1 _2776_/X sky130_fd_sc_hd__mux2_1
Xhold101 _1618_/X vssd1 vssd1 vccd1 vccd1 _3638_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1727_ _1727_/A _1727_/B vssd1 vssd1 vccd1 vccd1 _1739_/A sky130_fd_sc_hd__nand2_1
Xhold123 input20/X vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold134 _2732_/X vssd1 vssd1 vccd1 vccd1 _3263_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 _1656_/B vssd1 vssd1 vccd1 vccd1 _1667_/A sky130_fd_sc_hd__dlygate4sd3_1
X_1658_ input7/X hold33/X input9/X vssd1 vssd1 vccd1 vccd1 _1674_/C sky130_fd_sc_hd__and3_1
Xhold167 _3265_/Q vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _3310_/Q vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 _2764_/X vssd1 vssd1 vccd1 vccd1 _3292_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 _2748_/X vssd1 vssd1 vccd1 vccd1 _3278_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 _3608_/Q vssd1 vssd1 vccd1 vccd1 _1573_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3328_ _3333_/CLK _3328_/D vssd1 vssd1 vccd1 vccd1 _3328_/Q sky130_fd_sc_hd__dfxtp_1
X_1589_ _1589_/A vssd1 vssd1 vccd1 vccd1 _2130_/A sky130_fd_sc_hd__inv_2
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ _3521_/CLK _3259_/D vssd1 vssd1 vccd1 vccd1 _3259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2536__B1_N hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold690 _3411_/Q vssd1 vssd1 vccd1 vccd1 hold690/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1680__A1 hold45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2630_ _2360_/B hold606/X _2633_/S vssd1 vssd1 vccd1 vccd1 _2630_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2561_ _2574_/A _2561_/B vssd1 vssd1 vccd1 vccd1 _2561_/X sky130_fd_sc_hd__and2_2
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2492_ hold83/A _2510_/B _2489_/X _2491_/X vssd1 vssd1 vccd1 vccd1 _2492_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3113_ _3129_/A vssd1 vssd1 vccd1 vccd1 _3113_/Y sky130_fd_sc_hd__inv_2
X_3044_ _3049_/A vssd1 vssd1 vccd1 vccd1 _3044_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2844__S _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2620__A0 _2360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2828_ hold488/X _2355_/B _2829_/S vssd1 vssd1 vccd1 vccd1 _2828_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2759_ hold42/X hold30/X _2759_/S vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__mux2_1
XFILLER_0_5_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2687__A0 _2406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1662__A1 _2401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2611__A0 _2355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout73 _2087_/Y vssd1 vssd1 vccd1 vccd1 _2098_/S sky130_fd_sc_hd__buf_4
Xfanout95 hold820/X vssd1 vssd1 vccd1 vccd1 _2195_/A1 sky130_fd_sc_hd__buf_4
Xfanout84 _2532_/S1 vssd1 vssd1 vccd1 vccd1 _1912_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1653__A1 _2399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1992_ hold305/X hold303/X hold439/X hold312/X _2045_/S0 _2045_/S1 vssd1 vssd1 vccd1
+ vccd1 _1992_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_35_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3573_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2613_ _3519_/Q _2613_/B _3520_/Q vssd1 vssd1 vccd1 vccd1 _2881_/B sky130_fd_sc_hd__and3b_4
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3593_ _3607_/CLK _3593_/D _3084_/Y vssd1 vssd1 vccd1 vccd1 _3593_/Q sky130_fd_sc_hd__dfrtp_1
X_2544_ _3411_/Q _3402_/Q _3393_/Q _3438_/Q _1944_/B _1943_/A vssd1 vssd1 vccd1 vccd1
+ _2544_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_23_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2475_ _3610_/Q _2435_/A _2473_/X _2474_/X _2420_/X vssd1 vssd1 vccd1 vccd1 _2475_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2516__S0 _2532_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3027_ _3032_/A vssd1 vssd1 vccd1 vccd1 _3027_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2841__A0 _2358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2749__S _2749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2832__A0 _2098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1635__A1 hold45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2260_ _2363_/A _2259_/X _2228_/B vssd1 vssd1 vccd1 vccd1 _2270_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_20_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2191_ _2191_/A _2191_/B vssd1 vssd1 vccd1 vccd1 _2243_/B sky130_fd_sc_hd__or2_1
XFILLER_0_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1975_ _2315_/A1 _1975_/B vssd1 vssd1 vccd1 vccd1 _1975_/X sky130_fd_sc_hd__and2b_1
XANTENNA__2051__A1 _2036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout107_A hold117/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3576_ _3576_/CLK _3576_/D vssd1 vssd1 vccd1 vccd1 _3576_/Q sky130_fd_sc_hd__dfxtp_1
X_2527_ _2574_/A _2521_/X _2526_/X vssd1 vssd1 vccd1 vccd1 _2527_/X sky130_fd_sc_hd__o21a_1
X_2458_ _3609_/Q _2435_/A _2456_/X _2457_/X _2420_/X vssd1 vssd1 vccd1 vccd1 _2458_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__buf_4
Xhold49 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 input3/A sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ _1816_/B _1773_/Y _2384_/Y _1811_/S vssd1 vssd1 vccd1 vccd1 _3151_/D sky130_fd_sc_hd__a2bb2o_1
XANTENNA__1960__S1 _2045_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1760_ _1757_/B _2387_/C _1759_/X vssd1 vssd1 vccd1 vccd1 _1760_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_25_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold508 _3361_/Q vssd1 vssd1 vccd1 vccd1 hold508/X sky130_fd_sc_hd__dlygate4sd3_1
X_1691_ _1702_/A _1702_/B vssd1 vssd1 vccd1 vccd1 _1700_/B sky130_fd_sc_hd__or2_1
XFILLER_0_52_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold519 _2894_/X vssd1 vssd1 vccd1 vccd1 _3423_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3430_ _3438_/CLK _3430_/D vssd1 vssd1 vccd1 vccd1 _3430_/Q sky130_fd_sc_hd__dfxtp_1
X_3361_ _3516_/CLK _3361_/D vssd1 vssd1 vccd1 vccd1 _3361_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2312_ _3622_/Q _2070_/A _2121_/A _3623_/Q vssd1 vssd1 vccd1 vccd1 _2312_/X sky130_fd_sc_hd__a31o_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ _3332_/CLK _3292_/D vssd1 vssd1 vccd1 vccd1 _3292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2243_ _2729_/B _2243_/B vssd1 vssd1 vccd1 vccd1 _2243_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_79_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2174_ _2677_/B hold36/X vssd1 vssd1 vccd1 vccd1 _2578_/B sky130_fd_sc_hd__and2_2
XFILLER_0_73_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_50_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3433_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1958_ _2144_/C _3347_/Q _1956_/Y _2375_/A vssd1 vssd1 vccd1 vccd1 _2055_/S sky130_fd_sc_hd__o211a_4
X_1889_ _1923_/A _2363_/A vssd1 vssd1 vccd1 vccd1 _2613_/B sky130_fd_sc_hd__and2b_2
X_3628_ _3633_/CLK _3628_/D _3119_/Y vssd1 vssd1 vccd1 vccd1 _3628_/Q sky130_fd_sc_hd__dfstp_1
Xoutput39 _3439_/Q vssd1 vssd1 vccd1 vccd1 uart_tx sky130_fd_sc_hd__buf_12
X_3559_ _3559_/CLK _3559_/D _3053_/Y vssd1 vssd1 vccd1 vccd1 _3559_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2762__S _2769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2930_ _3090_/A vssd1 vssd1 vccd1 vccd1 _2930_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_84_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2861_ _2891_/A _2901_/B vssd1 vssd1 vccd1 vccd1 _2870_/S sky130_fd_sc_hd__and2_4
X_2792_ hold135/X _2802_/A1 _2799_/S vssd1 vssd1 vccd1 vccd1 _2792_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1812_ _2383_/A _1813_/B vssd1 vssd1 vccd1 vccd1 _1818_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_25_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1743_ _1886_/A _2383_/A _1886_/B vssd1 vssd1 vccd1 vccd1 _1743_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_7_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1674_ hold62/X _1674_/B _1674_/C vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__and3_4
XFILLER_0_40_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold305 _3222_/Q vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 _3237_/Q vssd1 vssd1 vccd1 vccd1 hold316/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 _3309_/Q vssd1 vssd1 vccd1 vccd1 hold327/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 _3279_/Q vssd1 vssd1 vccd1 vccd1 hold349/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 hold338/A vssd1 vssd1 vccd1 vccd1 hold338/X sky130_fd_sc_hd__buf_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3413_ _3413_/CLK _3413_/D vssd1 vssd1 vccd1 vccd1 _3413_/Q sky130_fd_sc_hd__dfxtp_1
X_3344_ _3610_/CLK _3344_/D _2919_/Y vssd1 vssd1 vccd1 vccd1 _3344_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 hold1052/X vssd1 vssd1 vccd1 vccd1 _1845_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2847__S _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _3320_/CLK _3275_/D vssd1 vssd1 vccd1 vccd1 _3275_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1016 _3519_/Q vssd1 vssd1 vccd1 vccd1 _1904_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1027 _3272_/Q vssd1 vssd1 vccd1 vccd1 _2742_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_2226_ _2208_/B _2223_/X _2224_/Y _2225_/X hold459/X vssd1 vssd1 vccd1 vccd1 _2226_/X
+ sky130_fd_sc_hd__a41o_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1049 _3443_/Q vssd1 vssd1 vccd1 vccd1 hold173/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2157_ _2157_/A _2157_/B vssd1 vssd1 vccd1 vccd1 _2157_/Y sky130_fd_sc_hd__nor2_1
X_2088_ _2077_/Y _2084_/Y _2092_/A vssd1 vssd1 vccd1 vccd1 _2088_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2582__S _2589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold850 _3499_/Q vssd1 vssd1 vccd1 vccd1 _2126_/A sky130_fd_sc_hd__buf_1
Xhold861 _2331_/X vssd1 vssd1 vccd1 vccd1 _3384_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 _2912_/X vssd1 vssd1 vccd1 vccd1 _3576_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout87_A _2532_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold894 _1701_/Y vssd1 vssd1 vccd1 vccd1 _3572_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 _2354_/X vssd1 vssd1 vccd1 vccd1 _3344_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2539__A2 hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3060_ _3061_/A vssd1 vssd1 vccd1 vccd1 _3060_/Y sky130_fd_sc_hd__inv_2
X_2011_ _2144_/C _2009_/X _2010_/Y vssd1 vssd1 vccd1 vccd1 _2011_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2913_ _3129_/A vssd1 vssd1 vccd1 vccd1 _2913_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_45_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2844_ _2105_/A hold552/X _2849_/S vssd1 vssd1 vccd1 vccd1 _2844_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2775_ hold307/X _2805_/A1 _2779_/S vssd1 vssd1 vccd1 vccd1 _2775_/X sky130_fd_sc_hd__mux2_1
Xhold124 _1672_/X vssd1 vssd1 vccd1 vccd1 _3603_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _3317_/Q vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__dlygate4sd3_1
X_1726_ _1839_/A _1726_/B vssd1 vssd1 vccd1 vccd1 _1727_/B sky130_fd_sc_hd__xnor2_1
Xhold102 hold102/A vssd1 vssd1 vccd1 vccd1 _2387_/A sky130_fd_sc_hd__buf_1
Xhold113 _2437_/A vssd1 vssd1 vccd1 vccd1 _1668_/B sky130_fd_sc_hd__dlygate4sd3_1
X_1657_ _1657_/A input4/X _1657_/C input6/X vssd1 vssd1 vccd1 vccd1 _1674_/B sky130_fd_sc_hd__and4_1
Xhold168 _2734_/X vssd1 vssd1 vccd1 vccd1 _3265_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 _2784_/X vssd1 vssd1 vccd1 vccd1 _3310_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 _3247_/Q vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
X_1588_ _1588_/A vssd1 vssd1 vccd1 vccd1 _1588_/Y sky130_fd_sc_hd__inv_2
Xhold179 _3254_/Q vssd1 vssd1 vccd1 vccd1 hold179/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3327_ _3504_/CLK _3327_/D vssd1 vssd1 vccd1 vccd1 _3327_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _3326_/CLK _3258_/D vssd1 vssd1 vccd1 vccd1 _3258_/Q sky130_fd_sc_hd__dfxtp_1
X_2209_ _2210_/C _2210_/B _2208_/Y vssd1 vssd1 vccd1 vccd1 _2209_/X sky130_fd_sc_hd__a21bo_1
X_3189_ _3433_/CLK _3189_/D vssd1 vssd1 vccd1 vccd1 _3189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold680 _3188_/Q vssd1 vssd1 vccd1 vccd1 hold680/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold691 _2880_/X vssd1 vssd1 vccd1 vccd1 _3411_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2560_ _3450_/Q _2510_/B _2557_/X _2559_/X vssd1 vssd1 vccd1 vccd1 _2561_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_50_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2491_ _3638_/Q _2510_/A _1643_/Y _3615_/Q _2490_/Y vssd1 vssd1 vccd1 vccd1 _2491_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2696__A1 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3112_ _3112_/A vssd1 vssd1 vccd1 vccd1 _3112_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_65_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3043_ _3049_/A vssd1 vssd1 vccd1 vccd1 _3043_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_85_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2827_ hold500/X _2357_/B _2829_/S vssd1 vssd1 vccd1 vccd1 _2827_/X sky130_fd_sc_hd__mux2_1
X_2758_ hold200/X _2808_/A1 _2759_/S vssd1 vssd1 vccd1 vccd1 _2758_/X sky130_fd_sc_hd__mux2_1
X_1709_ hold73/A _1871_/A vssd1 vssd1 vccd1 vccd1 _1709_/X sky130_fd_sc_hd__and2b_1
X_2689_ hold253/X _2801_/A1 _2697_/S vssd1 vssd1 vccd1 vccd1 _2689_/X sky130_fd_sc_hd__mux2_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_5_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3504_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_64_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout74 _2103_/Y vssd1 vssd1 vccd1 vccd1 _2104_/B sky130_fd_sc_hd__buf_4
Xfanout85 _3516_/Q vssd1 vssd1 vccd1 vccd1 _2532_/S1 sky130_fd_sc_hd__buf_4
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout96 _3483_/Q vssd1 vssd1 vccd1 vccd1 _2045_/S0 sky130_fd_sc_hd__buf_8
XFILLER_0_19_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1991_ hold376/X hold447/X hold392/X hold394/X _2045_/S0 _2045_/S1 vssd1 vssd1 vccd1
+ vccd1 _1991_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3592_ _3594_/CLK _3592_/D _3083_/Y vssd1 vssd1 vccd1 vccd1 _3592_/Q sky130_fd_sc_hd__dfrtp_1
X_2612_ _2356_/B hold628/X _2612_/S vssd1 vssd1 vccd1 vccd1 _2612_/X sky130_fd_sc_hd__mux2_1
X_2543_ _2542_/X _2541_/X _2546_/S vssd1 vssd1 vccd1 vccd1 _2543_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2474_ _3482_/Q _2507_/B _2508_/A vssd1 vssd1 vccd1 vccd1 _2474_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2669__A1 _2802_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3026_ _3032_/A vssd1 vssd1 vccd1 vccd1 _3026_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2516__S1 _2532_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2228__A_N _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2765__S _2769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1889__B _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2596__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2190_ _2219_/A _2221_/B _2222_/A vssd1 vssd1 vccd1 vccd1 _2191_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2823__A1 _2109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1974_ _1973_/X _1972_/X _2222_/A vssd1 vssd1 vccd1 vccd1 _1975_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3575_ _3575_/CLK _3575_/D _3069_/Y vssd1 vssd1 vccd1 vccd1 _3575_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2526_ hold89/A _2510_/B _2525_/X vssd1 vssd1 vccd1 vccd1 _2526_/X sky130_fd_sc_hd__a21o_1
X_2457_ _3481_/Q _2507_/B _2508_/A vssd1 vssd1 vccd1 vccd1 _2457_/X sky130_fd_sc_hd__o21a_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2585__S _2589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2388_ _1808_/A _1769_/B _2387_/X vssd1 vssd1 vccd1 vccd1 _2388_/X sky130_fd_sc_hd__a21o_1
XANTENNA__2814__A1 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3009_ _3110_/A vssd1 vssd1 vccd1 vccd1 _3009_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_66_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2805__A1 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold509 _2829_/X vssd1 vssd1 vccd1 vccd1 _3361_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1690_ _1704_/A _1704_/B vssd1 vssd1 vccd1 vccd1 _1702_/B sky130_fd_sc_hd__or2_1
XFILLER_0_52_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3360_ _3429_/CLK _3360_/D vssd1 vssd1 vccd1 vccd1 _3360_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2741__A0 _2801_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2311_ _1564_/Y _1977_/A _1988_/A vssd1 vssd1 vccd1 vccd1 _2314_/A sky130_fd_sc_hd__o21ai_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _3318_/CLK _3291_/D vssd1 vssd1 vccd1 vccd1 _3291_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2242_ _2223_/A _2242_/B _2242_/C _2242_/D vssd1 vssd1 vccd1 vccd1 _2242_/X sky130_fd_sc_hd__and4b_1
X_2173_ _2729_/B hold36/X _2172_/Y _2177_/A vssd1 vssd1 vccd1 vccd1 _2173_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1957_ _1957_/A _1957_/B vssd1 vssd1 vccd1 vccd1 _2375_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1888_ _1888_/A _1888_/B _1950_/C _1888_/D vssd1 vssd1 vccd1 vccd1 _2363_/A sky130_fd_sc_hd__and4_4
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3627_ _3627_/CLK hold46/X _3118_/Y vssd1 vssd1 vccd1 vccd1 _3627_/Q sky130_fd_sc_hd__dfrtp_2
X_3558_ _3559_/CLK _3558_/D _3052_/Y vssd1 vssd1 vccd1 vccd1 _3558_/Q sky130_fd_sc_hd__dfstp_1
X_2509_ _3585_/Q _2558_/B vssd1 vssd1 vccd1 vccd1 _2509_/X sky130_fd_sc_hd__or2_1
X_3489_ _3504_/CLK _3489_/D _2983_/Y vssd1 vssd1 vccd1 vccd1 _3489_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2723__A0 _2804_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_84_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2860_ _2356_/B hold694/X _2860_/S vssd1 vssd1 vccd1 vccd1 _2860_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1811_ _1810_/A _2383_/B _1811_/S vssd1 vssd1 vccd1 vccd1 _1813_/B sky130_fd_sc_hd__mux2_1
X_2791_ hold265/X _2801_/A1 _2799_/S vssd1 vssd1 vccd1 vccd1 _2791_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1742_ _1772_/B _1742_/B _1818_/A vssd1 vssd1 vccd1 vccd1 _1886_/B sky130_fd_sc_hd__nand3_2
Xhold306 _2684_/X vssd1 vssd1 vccd1 vccd1 _3222_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 _2701_/X vssd1 vssd1 vccd1 vccd1 _3237_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1673_ hold19/X hold9/X vssd1 vssd1 vccd1 vccd1 _2421_/B sky130_fd_sc_hd__nor2_4
Xhold339 _3282_/Q vssd1 vssd1 vccd1 vccd1 hold339/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 _2783_/X vssd1 vssd1 vccd1 vccd1 _3309_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3412_ _3516_/CLK _3412_/D vssd1 vssd1 vccd1 vccd1 _3412_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2714__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2190__A1 _2219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _3635_/CLK _3343_/D _2918_/Y vssd1 vssd1 vccd1 vccd1 _3343_/Q sky130_fd_sc_hd__dfrtp_1
Xhold1006 _3537_/Q vssd1 vssd1 vccd1 vccd1 _1853_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _3332_/CLK _3274_/D vssd1 vssd1 vccd1 vccd1 _3274_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1017 _3523_/Q vssd1 vssd1 vccd1 vccd1 _1587_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1028 _3552_/Q vssd1 vssd1 vccd1 vccd1 _1806_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_2225_ _2225_/A _2225_/B vssd1 vssd1 vccd1 vccd1 _2225_/X sky130_fd_sc_hd__or2_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2156_ _2155_/X _2129_/A _2158_/S vssd1 vssd1 vccd1 vccd1 _2156_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2863__S _2870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2087_ _2090_/A _2079_/X _2086_/X vssd1 vssd1 vccd1 vccd1 _2087_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2989_ _3054_/A vssd1 vssd1 vccd1 vccd1 _2989_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold862 _3469_/Q vssd1 vssd1 vccd1 vccd1 hold862/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2705__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold851 _2136_/X vssd1 vssd1 vccd1 vccd1 _3499_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 _3495_/Q vssd1 vssd1 vccd1 vccd1 _1589_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold840 _3580_/Q vssd1 vssd1 vccd1 vccd1 hold840/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 _3571_/Q vssd1 vssd1 vccd1 vccd1 _1702_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold895 _3570_/Q vssd1 vssd1 vccd1 vccd1 _1704_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2773__S _2779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_22_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2010_ _2010_/A _2144_/C vssd1 vssd1 vccd1 vccd1 _2010_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_29_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3635_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2912_ _1811_/S _1605_/Y _2911_/Y hold871/X vssd1 vssd1 vccd1 vccd1 _2912_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_85_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2843_ _2108_/Y hold704/X _2849_/S vssd1 vssd1 vccd1 vccd1 _2843_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2774_ hold161/X _2804_/A1 _2779_/S vssd1 vssd1 vccd1 vccd1 _2774_/X sky130_fd_sc_hd__mux2_1
X_1725_ _1843_/A hold84/X vssd1 vssd1 vccd1 vccd1 _1727_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold103 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 input14/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 hold125/A vssd1 vssd1 vccd1 vccd1 input27/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 _1668_/Y vssd1 vssd1 vccd1 vccd1 _1672_/S sky130_fd_sc_hd__clkbuf_2
Xhold136 _2792_/X vssd1 vssd1 vccd1 vccd1 _3317_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1656_ hold19/X _1656_/B vssd1 vssd1 vccd1 vccd1 _2165_/B sky130_fd_sc_hd__nor2_2
Xhold158 _2713_/X vssd1 vssd1 vccd1 vccd1 _3247_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _3593_/Q vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
X_1587_ _1587_/A vssd1 vssd1 vccd1 vccd1 _1885_/S sky130_fd_sc_hd__inv_2
Xhold169 _3319_/Q vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _3326_/CLK _3326_/D vssd1 vssd1 vccd1 vccd1 _3326_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _3326_/CLK _3257_/D vssd1 vssd1 vccd1 vccd1 _3257_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2208_ _2208_/A _2208_/B vssd1 vssd1 vccd1 vccd1 _2208_/Y sky130_fd_sc_hd__xnor2_1
X_3188_ _3431_/CLK _3188_/D vssd1 vssd1 vccd1 vccd1 _3188_/Q sky130_fd_sc_hd__dfxtp_1
X_2139_ _2139_/A _2139_/B vssd1 vssd1 vccd1 vccd1 _2143_/A sky130_fd_sc_hd__and2_1
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2768__S _2769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold681 _2642_/X vssd1 vssd1 vccd1 vccd1 _3188_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold670 _3171_/Q vssd1 vssd1 vccd1 vccd1 hold670/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 _3404_/Q vssd1 vssd1 vccd1 vccd1 hold692/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2490_ _2490_/A hold11/A vssd1 vssd1 vccd1 vccd1 _2490_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_49_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3111_ _3129_/A vssd1 vssd1 vccd1 vccd1 _3111_/Y sky130_fd_sc_hd__inv_2
X_3042_ _3054_/A vssd1 vssd1 vccd1 vccd1 _3042_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2826_ hold556/X _2360_/B _2829_/S vssd1 vssd1 vccd1 vccd1 _2826_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2908__A0 _2357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2757_ hold366/X _2807_/A1 _2759_/S vssd1 vssd1 vccd1 vccd1 _2757_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1708_ _1767_/S _1708_/B vssd1 vssd1 vccd1 vccd1 _1708_/X sky130_fd_sc_hd__xor2_1
X_2688_ _2800_/A _2719_/A vssd1 vssd1 vccd1 vccd1 _2697_/S sky130_fd_sc_hd__nor2_4
X_1639_ _2058_/D _2401_/A hold12/X vssd1 vssd1 vccd1 vccd1 _3623_/D sky130_fd_sc_hd__mux2_1
XANTENNA__2588__S _2589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ _3318_/CLK _3309_/D vssd1 vssd1 vccd1 vccd1 _3309_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout97 _3483_/Q vssd1 vssd1 vccd1 vccd1 _2221_/B sky130_fd_sc_hd__buf_6
XFILLER_0_24_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout86 _2532_/S0 vssd1 vssd1 vccd1 vccd1 _1944_/B sky130_fd_sc_hd__buf_8
Xfanout75 _2073_/X vssd1 vssd1 vccd1 vccd1 _2355_/B sky130_fd_sc_hd__buf_4
XFILLER_0_51_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1981__S0 _2045_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1990_ hold790/X _1989_/X _2055_/S vssd1 vssd1 vccd1 vccd1 _1990_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2611_ _2355_/B hold756/X _2612_/S vssd1 vssd1 vccd1 vccd1 _2611_/X sky130_fd_sc_hd__mux2_1
X_3591_ _3607_/CLK _3591_/D _3082_/Y vssd1 vssd1 vccd1 vccd1 _3591_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2542_ _3180_/Q _3429_/Q _3420_/Q _3162_/Q _1918_/B _1912_/B vssd1 vssd1 vccd1 vccd1
+ _2542_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_50_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1606__A _1607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2473_ _3606_/Q _2437_/A _2472_/X vssd1 vssd1 vccd1 vccd1 _2473_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_44_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3614_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1972__S0 _2221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3025_ _3032_/A vssd1 vssd1 vccd1 vccd1 _3025_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2809_ hold413/X _2406_/A _2809_/S vssd1 vssd1 vccd1 vccd1 _2809_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2781__S hold38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output43_A _2564_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2691__S _2697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1973_ _3251_/Q _3323_/Q _3314_/Q _3305_/Q _2049_/S0 _2195_/A1 vssd1 vssd1 vccd1
+ vccd1 _1973_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_7_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2587__A1 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3574_ _3574_/CLK _3574_/D _3068_/Y vssd1 vssd1 vccd1 vccd1 _3574_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2525_ hold99/A hold11/A _2522_/X _2524_/X _2559_/B vssd1 vssd1 vccd1 vccd1 _2525_/X
+ sky130_fd_sc_hd__o221a_1
X_2456_ _3605_/Q _2437_/A _2455_/X vssd1 vssd1 vccd1 vccd1 _2456_/X sky130_fd_sc_hd__a21o_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2866__S _2870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold29 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
X_2387_ _2387_/A _3149_/Q _2387_/C vssd1 vssd1 vccd1 vccd1 _2387_/X sky130_fd_sc_hd__and3_1
X_3008_ _3101_/A vssd1 vssd1 vccd1 vccd1 _3008_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2776__S _2779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1712__A_N _3454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2310_ _2310_/A _2310_/B vssd1 vssd1 vccd1 vccd1 _2324_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3290_ _3322_/CLK _3290_/D vssd1 vssd1 vccd1 vccd1 _3290_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2241_ _2708_/A _2241_/B vssd1 vssd1 vccd1 vccd1 _2242_/D sky130_fd_sc_hd__nand2_1
X_2172_ hold36/X _2222_/B vssd1 vssd1 vccd1 vccd1 _2172_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1956_ _2144_/C _2372_/S vssd1 vssd1 vccd1 vccd1 _1956_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_28_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1887_ _2490_/A _1808_/A _2911_/B vssd1 vssd1 vccd1 vccd1 _1888_/D sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout112_A hold123/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3626_ _3638_/CLK _3626_/D _3117_/Y vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__dfrtp_1
X_3557_ _3576_/CLK _3557_/D _3051_/Y vssd1 vssd1 vccd1 vccd1 _3557_/Q sky130_fd_sc_hd__dfstp_1
X_2508_ _2508_/A _2508_/B _2508_/C vssd1 vssd1 vccd1 vccd1 _2572_/C sky130_fd_sc_hd__and3_2
XANTENNA__2732__A1 _2802_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3488_ _3504_/CLK _3488_/D _2982_/Y vssd1 vssd1 vccd1 vccd1 _3488_/Q sky130_fd_sc_hd__dfrtp_4
X_2439_ _2436_/X _2508_/B _2438_/X _2437_/A _3604_/Q vssd1 vssd1 vccd1 vccd1 _2439_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2799__A1 hold30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2487__B1 _2479_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1810_ _1810_/A vssd1 vssd1 vccd1 vccd1 _1810_/Y sky130_fd_sc_hd__inv_2
X_2790_ _2790_/A _2790_/B vssd1 vssd1 vccd1 vccd1 _2799_/S sky130_fd_sc_hd__nor2_4
XFILLER_0_13_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1741_ _1888_/A _2228_/B vssd1 vssd1 vccd1 vccd1 _2383_/A sky130_fd_sc_hd__nand2_2
X_1672_ _2576_/A _3603_/Q _1672_/S vssd1 vssd1 vccd1 vccd1 _1672_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold307 _3302_/Q vssd1 vssd1 vccd1 vccd1 hold307/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 _3448_/Q vssd1 vssd1 vccd1 vccd1 _1730_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3411_ _3432_/CLK _3411_/D vssd1 vssd1 vccd1 vccd1 _3411_/Q sky130_fd_sc_hd__dfxtp_1
Xhold318 _3611_/Q vssd1 vssd1 vccd1 vccd1 _2358_/A sky130_fd_sc_hd__dlygate4sd3_1
X_3342_ _3432_/CLK _3342_/D vssd1 vssd1 vccd1 vccd1 _3342_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2190__A2 _2221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _3318_/CLK _3273_/D vssd1 vssd1 vccd1 vccd1 _3273_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1007 _3498_/Q vssd1 vssd1 vccd1 vccd1 _2119_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 _3577_/Q vssd1 vssd1 vccd1 vccd1 hold1018/X sky130_fd_sc_hd__dlygate4sd3_1
X_2224_ _2225_/A _2225_/B vssd1 vssd1 vccd1 vccd1 _2224_/Y sky130_fd_sc_hd__nand2_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1029 _3500_/Q vssd1 vssd1 vccd1 vccd1 _2335_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2155_ _2155_/A _2155_/B _2155_/C vssd1 vssd1 vccd1 vccd1 _2155_/X sky130_fd_sc_hd__and3_1
XFILLER_0_88_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2086_ _2064_/B _2085_/X _2082_/X _2067_/B vssd1 vssd1 vccd1 vccd1 _2086_/X sky130_fd_sc_hd__a211o_1
XANTENNA__2650__A0 _2104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2164__B _3577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2988_ _3127_/A vssd1 vssd1 vccd1 vccd1 _2988_/Y sky130_fd_sc_hd__inv_2
X_1939_ _3511_/Q _1939_/B vssd1 vssd1 vccd1 vccd1 _1939_/X sky130_fd_sc_hd__or2_1
Xhold830 _1697_/Y vssd1 vssd1 vccd1 vccd1 _3462_/D sky130_fd_sc_hd__clkbuf_2
X_3609_ _3610_/CLK _3609_/D _3100_/Y vssd1 vssd1 vccd1 vccd1 _3609_/Q sky130_fd_sc_hd__dfrtp_1
Xhold841 _1688_/X vssd1 vssd1 vccd1 vccd1 _3590_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold863 _2252_/X vssd1 vssd1 vccd1 vccd1 _3469_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold852 _3466_/Q vssd1 vssd1 vccd1 vccd1 hold852/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 _1704_/Y vssd1 vssd1 vccd1 vccd1 hold896/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 _1702_/Y vssd1 vssd1 vccd1 vccd1 hold885/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 _2151_/Y vssd1 vssd1 vccd1 vccd1 _3495_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2641__A0 _2357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2880__A0 _2356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1683__A1 hold75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2632__A0 _2355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2911_ _3054_/A _2911_/B _2911_/C vssd1 vssd1 vccd1 vccd1 _2911_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_45_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2842_ _2087_/Y hold640/X _2849_/S vssd1 vssd1 vccd1 vccd1 _2842_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2773_ hold336/X _2803_/A1 _2779_/S vssd1 vssd1 vccd1 vccd1 _2773_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3096__A _3124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1724_ _3524_/Q _1724_/B vssd1 vssd1 vccd1 vccd1 _1724_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1609__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold104 _1612_/A vssd1 vssd1 vccd1 vccd1 _1624_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 input27/X vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_hold50_A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold115 _1671_/X vssd1 vssd1 vccd1 vccd1 _3604_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 _3299_/Q vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__dlygate4sd3_1
X_1655_ hold92/X hold50/X _1655_/C hold8/X vssd1 vssd1 vccd1 vccd1 _1656_/B sky130_fd_sc_hd__or4b_1
Xhold159 _3274_/Q vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 _1686_/X vssd1 vssd1 vccd1 vccd1 _3593_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1586_ _1840_/A vssd1 vssd1 vccd1 vccd1 _1879_/A sky130_fd_sc_hd__inv_2
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2699__A0 _2801_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ _3330_/CLK _3325_/D vssd1 vssd1 vccd1 vccd1 _3325_/Q sky130_fd_sc_hd__dfxtp_1
X_3256_ _3326_/CLK _3256_/D vssd1 vssd1 vccd1 vccd1 _3256_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2207_ _2204_/A _2204_/B _2213_/B vssd1 vssd1 vccd1 vccd1 _2210_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__2874__S _2880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3187_ _3521_/CLK _3187_/D vssd1 vssd1 vccd1 vccd1 _3187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2138_ _2138_/A _2138_/B vssd1 vssd1 vccd1 vccd1 _3498_/D sky130_fd_sc_hd__and2_1
X_2069_ _2059_/Y _2068_/Y _2092_/A vssd1 vssd1 vccd1 vccd1 _2069_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2623__A0 _2356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold671 _2623_/X vssd1 vssd1 vccd1 vccd1 _3171_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold660 _3195_/Q vssd1 vssd1 vccd1 vccd1 hold660/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 _2873_/X vssd1 vssd1 vccd1 vccd1 _3404_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 _3385_/Q vssd1 vssd1 vccd1 vccd1 hold682/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2784__S hold38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1665__A1 _2576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3110_ _3110_/A vssd1 vssd1 vccd1 vccd1 _3110_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2528__S0 _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3041_ _3049_/A vssd1 vssd1 vccd1 vccd1 _3041_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2694__S _2697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2853__A0 _2098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2605__A0 _2098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2825_ hold610/X _2104_/B _2829_/S vssd1 vssd1 vccd1 vccd1 _2825_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2756_ hold282/X _2806_/A1 _2759_/S vssd1 vssd1 vccd1 vccd1 _2756_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2869__S _2870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1707_ _1704_/B _1706_/Y _3462_/D vssd1 vssd1 vccd1 vccd1 _3569_/D sky130_fd_sc_hd__a21oi_1
X_2687_ _2406_/A hold425/X _2687_/S vssd1 vssd1 vccd1 vccd1 _2687_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1638_ _2387_/A hold75/X hold12/X vssd1 vssd1 vccd1 vccd1 _3624_/D sky130_fd_sc_hd__mux2_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1569_ _1569_/A vssd1 vssd1 vccd1 vccd1 _1569_/Y sky130_fd_sc_hd__inv_2
X_3308_ _3319_/CLK _3308_/D vssd1 vssd1 vccd1 vccd1 _3308_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2519__S0 _1918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3239_ _3326_/CLK _3239_/D vssd1 vssd1 vccd1 vccd1 _3239_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2844__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1647__A1 hold45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout98 _3483_/Q vssd1 vssd1 vccd1 vccd1 _2049_/S0 sky130_fd_sc_hd__clkbuf_4
Xfanout87 _2532_/S0 vssd1 vssd1 vccd1 vccd1 _1918_/B sky130_fd_sc_hd__buf_6
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout76 _2072_/Y vssd1 vssd1 vccd1 vccd1 _2357_/B sky130_fd_sc_hd__buf_4
XANTENNA__2779__S _2779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold490 _3429_/Q vssd1 vssd1 vccd1 vccd1 hold490/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1981__S1 _2045_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2835__A0 _2104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1638__A1 hold75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3590_ _3590_/CLK _3590_/D _3081_/Y vssd1 vssd1 vccd1 vccd1 _3590_/Q sky130_fd_sc_hd__dfrtp_1
X_2610_ _2357_/B hold748/X _2612_/S vssd1 vssd1 vccd1 vccd1 _2610_/X sky130_fd_sc_hd__mux2_1
X_2541_ _3379_/Q _3361_/Q _3370_/Q _3198_/Q _1918_/B _1912_/B vssd1 vssd1 vccd1 vccd1
+ _2541_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2366__A2 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2689__S _2697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2472_ _3583_/Q _2558_/B _2508_/B _2471_/X vssd1 vssd1 vccd1 vccd1 _2472_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1606__B _1607_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1972__S1 _2195_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3024_ _3032_/A vssd1 vssd1 vccd1 vccd1 _3024_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_13_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3324_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2054__A1 _2144_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2808_ hold230/X _2808_/A1 _2809_/S vssd1 vssd1 vccd1 vccd1 _2808_/X sky130_fd_sc_hd__mux2_1
X_2739_ hold343/X _2406_/A _2739_/S vssd1 vssd1 vccd1 vccd1 _2739_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1963__S1 _2219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2363__A _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1972_ _3296_/Q _3287_/Q _3278_/Q _3269_/Q _2221_/B _2195_/A1 vssd1 vssd1 vccd1 vccd1
+ _1972_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_15_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3573_ _3573_/CLK _3573_/D _3067_/Y vssd1 vssd1 vccd1 vccd1 _3573_/Q sky130_fd_sc_hd__dfrtp_1
X_2524_ _3598_/Q _2438_/B _2572_/C _2523_/X vssd1 vssd1 vccd1 vccd1 _2524_/X sky130_fd_sc_hd__o211a_1
X_2455_ _3582_/Q _2558_/B _2508_/B _2454_/X vssd1 vssd1 vccd1 vccd1 _2455_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_11_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2386_ _2184_/A _1957_/B _2146_/A _2381_/X vssd1 vssd1 vccd1 vccd1 _2386_/X sky130_fd_sc_hd__a22o_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__buf_2
XFILLER_0_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2882__S _2890_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3007_ _3101_/A vssd1 vssd1 vccd1 vccd1 _3007_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_61_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1961__S _2036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2792__S _2799_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3652__A _3655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ _2240_/A _2240_/B vssd1 vssd1 vccd1 vccd1 _3473_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2171_ _2171_/A _2171_/B vssd1 vssd1 vccd1 vccd1 _2222_/B sky130_fd_sc_hd__or2_1
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1955_ _2381_/A _2381_/B _2381_/C _1955_/D vssd1 vssd1 vccd1 vccd1 _2372_/S sky130_fd_sc_hd__or4_2
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1886_ _1886_/A _1886_/B _1886_/C vssd1 vssd1 vccd1 vccd1 _2911_/B sky130_fd_sc_hd__or3_1
XFILLER_0_3_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3625_ _3627_/CLK _3625_/D _3116_/Y vssd1 vssd1 vccd1 vccd1 _3625_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout105_A hold75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3556_ _3576_/CLK _3556_/D _3050_/Y vssd1 vssd1 vccd1 vccd1 _3556_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__2877__S _2880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2507_ hold52/A _2507_/B _2507_/C vssd1 vssd1 vccd1 vccd1 _2508_/C sky130_fd_sc_hd__and3_1
X_3487_ _3504_/CLK _3487_/D _2981_/Y vssd1 vssd1 vccd1 vccd1 _3487_/Q sky130_fd_sc_hd__dfrtp_1
X_2438_ _3593_/Q _2438_/B vssd1 vssd1 vccd1 vccd1 _2438_/X sky130_fd_sc_hd__or2_1
X_2369_ _3627_/Q hold99/X hold72/X vssd1 vssd1 vccd1 vccd1 _2370_/A sky130_fd_sc_hd__or3_2
XFILLER_0_78_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2360__B _2360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2787__S hold38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2487__A1 _1908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3647__A _3655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1740_ _2381_/B _2381_/C vssd1 vssd1 vccd1 vccd1 _2228_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_80_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold308 _2775_/X vssd1 vssd1 vccd1 vccd1 _3302_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1671_ _2399_/A _3604_/Q _1672_/S vssd1 vssd1 vccd1 vccd1 _1671_/X sky130_fd_sc_hd__mux2_1
X_3410_ _3431_/CLK _3410_/D vssd1 vssd1 vccd1 vccd1 _3410_/Q sky130_fd_sc_hd__dfxtp_1
Xhold319 _3215_/Q vssd1 vssd1 vccd1 vccd1 hold319/X sky130_fd_sc_hd__dlygate4sd3_1
X_3341_ _3431_/CLK _3341_/D vssd1 vssd1 vccd1 vccd1 _3341_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2697__S _2697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _3319_/CLK _3272_/D vssd1 vssd1 vccd1 vccd1 _3272_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1008 _3538_/Q vssd1 vssd1 vccd1 vccd1 _1855_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1019 _3451_/Q vssd1 vssd1 vccd1 vccd1 _1716_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ _2223_/A _2242_/B _2242_/C _2223_/D vssd1 vssd1 vccd1 vccd1 _2223_/X sky130_fd_sc_hd__and4_1
X_2154_ _2158_/S _2152_/Y hold931/X vssd1 vssd1 vccd1 vccd1 _2154_/X sky130_fd_sc_hd__o21a_1
X_2085_ _2083_/Y _2084_/Y _2091_/S vssd1 vssd1 vccd1 vccd1 _2085_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2987_ _3054_/A vssd1 vssd1 vccd1 vccd1 _2987_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1938_ _1934_/B _1937_/Y _1929_/A _1935_/B vssd1 vssd1 vccd1 vccd1 _3513_/D sky130_fd_sc_hd__a2bb2o_1
X_1869_ _1583_/Y _1846_/Y _1837_/Y vssd1 vssd1 vccd1 vccd1 _1869_/X sky130_fd_sc_hd__a21o_1
Xhold820 _3484_/Q vssd1 vssd1 vccd1 vccd1 hold820/X sky130_fd_sc_hd__dlygate4sd3_1
X_3608_ _3610_/CLK _3608_/D _3099_/Y vssd1 vssd1 vccd1 vccd1 _3608_/Q sky130_fd_sc_hd__dfrtp_1
Xhold842 _3526_/Q vssd1 vssd1 vccd1 vccd1 _1840_/A sky130_fd_sc_hd__buf_1
Xhold853 _2254_/X vssd1 vssd1 vccd1 vccd1 _3467_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold831 _3555_/Q vssd1 vssd1 vccd1 vccd1 _1791_/A sky130_fd_sc_hd__buf_1
Xhold864 _3152_/Q vssd1 vssd1 vccd1 vccd1 _1808_/A sky130_fd_sc_hd__buf_1
X_3539_ _3575_/CLK _3539_/D _3033_/Y vssd1 vssd1 vccd1 vccd1 _3539_/Q sky130_fd_sc_hd__dfrtp_1
Xhold886 _1703_/Y vssd1 vssd1 vccd1 vccd1 _3571_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 _1705_/Y vssd1 vssd1 vccd1 vccd1 _3570_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 _3347_/Q vssd1 vssd1 vccd1 vccd1 _1957_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__2013__S0 _2045_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2355__B _2355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2004__S0 _2045_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2910_ _2356_/B hold616/X _2910_/S vssd1 vssd1 vccd1 vccd1 _2910_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2841_ _2358_/B hold696/X _2849_/S vssd1 vssd1 vccd1 vccd1 _2841_/X sky130_fd_sc_hd__mux2_1
X_2772_ hold137/X _2802_/A1 _2779_/S vssd1 vssd1 vccd1 vccd1 _2772_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1723_ _1865_/A _3450_/Q vssd1 vssd1 vccd1 vccd1 _1723_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_13_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_38_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3579_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1609__B input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold116 hold116/A vssd1 vssd1 vccd1 vccd1 input29/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 _1624_/X vssd1 vssd1 vccd1 vccd1 _1625_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _2772_/X vssd1 vssd1 vccd1 vccd1 _3299_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 input5/A sky130_fd_sc_hd__dlygate4sd3_1
X_1654_ _2358_/A _2576_/A hold53/X vssd1 vssd1 vccd1 vccd1 _3611_/D sky130_fd_sc_hd__mux2_1
Xhold127 _2742_/X vssd1 vssd1 vccd1 vccd1 _3272_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1585_ _1877_/A vssd1 vssd1 vccd1 vccd1 _1585_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3324_ _3324_/CLK hold48/X vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dfxtp_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3320_/CLK _3255_/D vssd1 vssd1 vccd1 vccd1 _3255_/Q sky130_fd_sc_hd__dfxtp_1
X_2206_ _2210_/C _2206_/B vssd1 vssd1 vccd1 vccd1 _2213_/B sky130_fd_sc_hd__and2_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _3408_/CLK _3186_/D vssd1 vssd1 vccd1 vccd1 _3186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2137_ _2119_/B _2139_/A _2139_/B _2119_/A vssd1 vssd1 vccd1 vccd1 _2138_/B sky130_fd_sc_hd__a31o_1
X_2068_ _3545_/Q _2084_/B vssd1 vssd1 vccd1 vccd1 _2068_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2890__S _2890_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold650 _3163_/Q vssd1 vssd1 vccd1 vccd1 hold650/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 _3185_/Q vssd1 vssd1 vccd1 vccd1 hold672/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 _2651_/X vssd1 vssd1 vccd1 vccd1 _3195_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 _3393_/Q vssd1 vssd1 vccd1 vccd1 hold694/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 _2852_/X vssd1 vssd1 vccd1 vccd1 _3385_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2862__A1 _2358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output66_A _2552_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2528__S1 _2532_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3040_ _3049_/A vssd1 vssd1 vccd1 vccd1 _3040_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_81_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2824_ hold496/X _2105_/A _2829_/S vssd1 vssd1 vccd1 vccd1 _2824_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2464__S0 _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2755_ hold314/X _2805_/A1 _2759_/S vssd1 vssd1 vccd1 vccd1 _2755_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1706_ _1689_/A _1708_/B _1689_/B vssd1 vssd1 vccd1 vccd1 _1706_/Y sky130_fd_sc_hd__o21ai_1
X_2686_ _2808_/A1 hold299/X _2687_/S vssd1 vssd1 vccd1 vccd1 _2686_/X sky130_fd_sc_hd__mux2_1
X_1637_ hold72/X hold70/X hold12/X vssd1 vssd1 vccd1 vccd1 _3625_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_1_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3307_ _3318_/CLK _3307_/D vssd1 vssd1 vccd1 vccd1 _3307_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2885__S _2890_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1568_ _1568_/A vssd1 vssd1 vccd1 vccd1 _1568_/Y sky130_fd_sc_hd__inv_2
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2519__S1 _2532_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3238_ _3326_/CLK _3238_/D vssd1 vssd1 vccd1 vccd1 _3238_/Q sky130_fd_sc_hd__dfxtp_1
X_3169_ _3432_/CLK _3169_/D vssd1 vssd1 vccd1 vccd1 _3169_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2285__D_N _1623_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout88 hold817/X vssd1 vssd1 vccd1 vccd1 _2532_/S0 sky130_fd_sc_hd__buf_6
Xfanout77 _2058_/X vssd1 vssd1 vccd1 vccd1 _2356_/B sky130_fd_sc_hd__buf_4
Xfanout99 hold940/X vssd1 vssd1 vccd1 vccd1 _2144_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold480 _3586_/Q vssd1 vssd1 vccd1 vccd1 _2338_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold491 _2900_/X vssd1 vssd1 vccd1 vccd1 _3429_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2795__S _2799_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2599__A0 _2357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3655__A _3655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2446__S0 _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2540_ _2574_/A _2534_/X _2535_/X _2539_/X vssd1 vssd1 vccd1 vccd1 _2540_/X sky130_fd_sc_hd__o22a_2
XFILLER_0_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2471_ _3595_/Q _2438_/B _2558_/C _3344_/Q vssd1 vssd1 vccd1 vccd1 _2471_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_76_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3023_ _3032_/A vssd1 vssd1 vccd1 vccd1 _3023_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2826__A1 _2360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2807_ hold415/X _2807_/A1 _2809_/S vssd1 vssd1 vccd1 vccd1 _2807_/X sky130_fd_sc_hd__mux2_1
X_2738_ hold202/X _2808_/A1 _2739_/S vssd1 vssd1 vccd1 vccd1 _2738_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2762__A0 _2802_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2669_ hold182/X _2802_/A1 _2676_/S vssd1 vssd1 vccd1 vccd1 _2669_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2817__A1 _2357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2428__S0 _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2808__A1 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2284__A2 _2270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1971_ _1969_/X _1970_/X _2036_/S vssd1 vssd1 vccd1 vccd1 _1971_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_36_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3572_ _3573_/CLK _3572_/D _3066_/Y vssd1 vssd1 vccd1 vccd1 _3572_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2523_ _3586_/Q _2558_/B _2558_/C _3380_/Q vssd1 vssd1 vccd1 vccd1 _2523_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_51_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2744__A0 _2804_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2454_ _3594_/Q _2438_/B _2558_/C _3345_/Q vssd1 vssd1 vccd1 vccd1 _2454_/X sky130_fd_sc_hd__o22a_1
X_2385_ _1811_/S _2911_/C _2385_/B1 vssd1 vssd1 vccd1 vccd1 _3148_/D sky130_fd_sc_hd__a21o_1
Xinput1 uart_rx vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3006_ _3101_/A vssd1 vssd1 vccd1 vccd1 _3006_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2183__B _2198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2358__B _2358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2726__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2170_ _3488_/Q _2677_/B _2729_/B vssd1 vssd1 vccd1 vccd1 _2171_/B sky130_fd_sc_hd__a21oi_1
X_1954_ _2130_/A _2152_/A vssd1 vssd1 vccd1 vccd1 _1955_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1885_ _1836_/A _1837_/A _1885_/S vssd1 vssd1 vccd1 vccd1 _3523_/D sky130_fd_sc_hd__mux2_1
X_3624_ _3638_/CLK _3624_/D _3115_/Y vssd1 vssd1 vccd1 vccd1 _3624_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2717__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3555_ _3555_/CLK _3555_/D _3049_/Y vssd1 vssd1 vccd1 vccd1 _3555_/Q sky130_fd_sc_hd__dfrtp_1
X_3486_ _3590_/CLK _3486_/D _2980_/Y vssd1 vssd1 vccd1 vccd1 _3486_/Q sky130_fd_sc_hd__dfrtp_1
X_2506_ hold84/A hold35/A hold20/A vssd1 vssd1 vccd1 vccd1 _2506_/X sky130_fd_sc_hd__and3_1
X_2437_ _2437_/A _2437_/B vssd1 vssd1 vccd1 vccd1 _2508_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2368_ _3343_/Q _2367_/X hold800/X vssd1 vssd1 vccd1 vccd1 _2368_/X sky130_fd_sc_hd__o21ba_1
X_2299_ hold89/X hold87/X hold22/X vssd1 vssd1 vccd1 vccd1 _3446_/D sky130_fd_sc_hd__mux2_1
XANTENNA__2893__S _2900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2270__C _2270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1670_ _2400_/A _3605_/Q _1672_/S vssd1 vssd1 vccd1 vccd1 _1670_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold309 _3268_/Q vssd1 vssd1 vccd1 vccd1 hold309/X sky130_fd_sc_hd__dlygate4sd3_1
X_3340_ _3432_/CLK _3340_/D vssd1 vssd1 vccd1 vccd1 _3340_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3321_/CLK _3271_/D vssd1 vssd1 vccd1 vccd1 _3271_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1009 _3554_/Q vssd1 vssd1 vccd1 vccd1 _1771_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _2222_/A _2222_/B vssd1 vssd1 vccd1 vccd1 _2223_/D sky130_fd_sc_hd__xor2_1
XFILLER_0_17_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2153_ _3493_/Q _3492_/Q _2375_/A _2148_/B _2130_/B vssd1 vssd1 vccd1 vccd1 _2153_/X
+ sky130_fd_sc_hd__a41o_1
X_2084_ _3543_/Q _2084_/B vssd1 vssd1 vccd1 vccd1 _2084_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2986_ _3054_/A vssd1 vssd1 vccd1 vccd1 _2986_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1937_ _1931_/A _1931_/B _1935_/Y vssd1 vssd1 vccd1 vccd1 _1937_/Y sky130_fd_sc_hd__o21ai_1
X_1868_ _1867_/Y _1865_/B _1848_/A _1836_/A vssd1 vssd1 vccd1 vccd1 _1868_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_31_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold821 _2195_/X vssd1 vssd1 vccd1 vccd1 _3484_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold810 _1903_/Y vssd1 vssd1 vccd1 vccd1 _3520_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2888__S _2890_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3607_ _3607_/CLK _3607_/D _3098_/Y vssd1 vssd1 vccd1 vccd1 _3607_/Q sky130_fd_sc_hd__dfrtp_1
X_3538_ _3632_/CLK _3538_/D _3032_/Y vssd1 vssd1 vccd1 vccd1 _3538_/Q sky130_fd_sc_hd__dfrtp_1
Xhold843 _1880_/X vssd1 vssd1 vccd1 vccd1 _3526_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold854 _3589_/Q vssd1 vssd1 vccd1 vccd1 hold854/X sky130_fd_sc_hd__dlygate4sd3_1
X_1799_ _1791_/A _1801_/A _1798_/X vssd1 vssd1 vccd1 vccd1 _1799_/X sky130_fd_sc_hd__a21o_1
Xhold832 _1799_/X vssd1 vssd1 vccd1 vccd1 _3555_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 _3463_/Q vssd1 vssd1 vccd1 vccd1 hold898/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 _2329_/X vssd1 vssd1 vccd1 vccd1 hold876/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 _2388_/X vssd1 vssd1 vccd1 vccd1 _3152_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 _3351_/Q vssd1 vssd1 vccd1 vccd1 _2144_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3469_ _3574_/CLK _3469_/D _2963_/Y vssd1 vssd1 vccd1 vccd1 _3469_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2013__S1 _2045_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_8_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3320_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2798__S _2799_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2004__S1 _2045_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2093__B1 _2064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2840_ _3520_/Q _3519_/Q _2871_/C _2830_/B vssd1 vssd1 vccd1 vccd1 _2849_/S sky130_fd_sc_hd__or4b_4
X_2771_ hold269/X _2801_/A1 _2779_/S vssd1 vssd1 vccd1 vccd1 _2771_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1722_ _1717_/B _1848_/A vssd1 vssd1 vccd1 vccd1 _1722_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold117 input29/X vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__clkbuf_2
X_1653_ _1570_/A _2399_/A hold53/X vssd1 vssd1 vccd1 vccd1 _3612_/D sky130_fd_sc_hd__mux2_1
Xhold106 _1626_/B vssd1 vssd1 vccd1 vccd1 _1666_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2501__S _2546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold139 _3623_/Q vssd1 vssd1 vccd1 vccd1 _2058_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold128 _3595_/Q vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
X_1584_ _1845_/A vssd1 vssd1 vccd1 vccd1 _1584_/Y sky130_fd_sc_hd__inv_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3323_ _3324_/CLK _3323_/D vssd1 vssd1 vccd1 vccd1 _3323_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ _3408_/CLK _3254_/D vssd1 vssd1 vccd1 vccd1 _3254_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _2205_/A _2205_/B vssd1 vssd1 vccd1 vccd1 _2206_/B sky130_fd_sc_hd__or2_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ _3433_/CLK _3185_/D vssd1 vssd1 vccd1 vccd1 _3185_/Q sky130_fd_sc_hd__dfxtp_1
X_2136_ _2126_/A _2138_/A _2135_/X vssd1 vssd1 vccd1 vccd1 _2136_/X sky130_fd_sc_hd__a21o_1
X_2067_ _2090_/A _2067_/B vssd1 vssd1 vccd1 vccd1 _2106_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_88_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_76_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2969_ _3061_/A vssd1 vssd1 vccd1 vccd1 _2969_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_4_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold651 _2615_/X vssd1 vssd1 vccd1 vccd1 _3163_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 _3170_/Q vssd1 vssd1 vccd1 vccd1 hold662/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold640 _3372_/Q vssd1 vssd1 vccd1 vccd1 hold640/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 _3405_/Q vssd1 vssd1 vccd1 vccd1 hold684/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 _2860_/X vssd1 vssd1 vccd1 vccd1 _3393_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 _2639_/X vssd1 vssd1 vccd1 vccd1 _3185_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1984__S0 _2221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2302__A1 _2401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2823_ hold520/X _2109_/B _2829_/S vssd1 vssd1 vccd1 vccd1 _2823_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2754_ hold165/X _2804_/A1 _2759_/S vssd1 vssd1 vccd1 vccd1 _2754_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_81_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2464__S1 _1943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1705_ _1702_/B hold896/X _3462_/D vssd1 vssd1 vccd1 vccd1 _1705_/Y sky130_fd_sc_hd__a21oi_1
X_2685_ _2807_/A1 hold411/X _2687_/S vssd1 vssd1 vccd1 vccd1 _2685_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1636_ hold99/X hold87/X hold12/X vssd1 vssd1 vccd1 vccd1 _3626_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_1_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1567_ _3615_/Q vssd1 vssd1 vccd1 vccd1 _1567_/Y sky130_fd_sc_hd__inv_2
X_3306_ _3324_/CLK hold41/X vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__dfxtp_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _3320_/CLK _3237_/D vssd1 vssd1 vccd1 vccd1 _3237_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3168_ _3438_/CLK _3168_/D vssd1 vssd1 vccd1 vccd1 _3168_/Q sky130_fd_sc_hd__dfxtp_1
X_2119_ _2119_/A _2119_/B _2139_/A vssd1 vssd1 vccd1 vccd1 _2135_/C sky130_fd_sc_hd__and3_1
X_3099_ _3101_/A vssd1 vssd1 vccd1 vccd1 _3099_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_71_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout78 hold10/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__buf_4
Xfanout89 _2225_/A vssd1 vssd1 vccd1 vccd1 _2315_/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_32_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold481 _2338_/Y vssd1 vssd1 vccd1 vccd1 _3380_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold470 _1909_/Y vssd1 vssd1 vccd1 vccd1 hold470/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 _3340_/Q vssd1 vssd1 vccd1 vccd1 hold492/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2446__S1 _1943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2771__A1 _2801_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2470_ _1908_/D _2469_/X _2462_/X vssd1 vssd1 vccd1 vccd1 _2470_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3022_ _3032_/A vssd1 vssd1 vccd1 vccd1 _3022_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_58_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout128_A _3057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2806_ hold312/X _2806_/A1 _2809_/S vssd1 vssd1 vccd1 vccd1 _2806_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_22_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3632_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2737_ hold309/X _2807_/A1 _2739_/S vssd1 vssd1 vccd1 vccd1 _2737_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2668_ hold292/X _2801_/A1 _2676_/S vssd1 vssd1 vccd1 vccd1 _2668_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2896__S _2900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1619_ _1768_/S _2401_/A _1622_/S vssd1 vssd1 vccd1 vccd1 _1619_/X sky130_fd_sc_hd__mux2_1
X_2599_ _2357_/B hold624/X _2601_/S vssd1 vssd1 vccd1 vccd1 _2599_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2514__A1 _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2428__S1 _1943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2753__A1 _2803_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1970_ hold299/X hold319/X hold212/X hold230/X _3483_/Q _2045_/S1 vssd1 vssd1 vccd1
+ vccd1 _1970_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_28_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2570__A _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3571_ _3571_/CLK _3571_/D _3065_/Y vssd1 vssd1 vccd1 vccd1 _3571_/Q sky130_fd_sc_hd__dfrtp_1
X_2522_ hold90/A _1643_/Y hold11/A vssd1 vssd1 vccd1 vccd1 _2522_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_51_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2453_ _1908_/D _2452_/X _2445_/X vssd1 vssd1 vccd1 vccd1 _2453_/X sky130_fd_sc_hd__a21o_1
X_2384_ _2911_/C vssd1 vssd1 vccd1 vccd1 _2384_/Y sky130_fd_sc_hd__inv_2
Xinput2 wb_rst_i vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_4
X_3005_ _3110_/A vssd1 vssd1 vccd1 vccd1 _3005_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2680__A0 _2802_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2735__A1 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output41_A _2434_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2662__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1953_ _2130_/A _2152_/A vssd1 vssd1 vccd1 vccd1 _2379_/C sky130_fd_sc_hd__and2_1
XFILLER_0_71_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1884_ _1837_/A _1838_/Y _1883_/X _1883_/A _1836_/A vssd1 vssd1 vccd1 vccd1 _1884_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__2504__S _3517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3623_ _3627_/CLK _3623_/D _3114_/Y vssd1 vssd1 vccd1 vccd1 _3623_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3554_ _3571_/CLK _3554_/D _3048_/Y vssd1 vssd1 vccd1 vccd1 _3554_/Q sky130_fd_sc_hd__dfrtp_1
X_3485_ _3605_/CLK _3485_/D _2979_/Y vssd1 vssd1 vccd1 vccd1 _3485_/Q sky130_fd_sc_hd__dfrtp_1
X_2505_ _2504_/X _2501_/X _3518_/Q vssd1 vssd1 vccd1 vccd1 _2505_/X sky130_fd_sc_hd__mux2_1
X_2436_ _3581_/Q _2558_/B _2558_/C _3384_/Q vssd1 vssd1 vccd1 vccd1 _2436_/X sky130_fd_sc_hd__o22a_1
X_2367_ _2362_/X _2367_/B _2367_/C _2367_/D vssd1 vssd1 vccd1 vccd1 _2367_/X sky130_fd_sc_hd__and4b_1
X_2298_ hold73/X hold45/X hold22/X vssd1 vssd1 vccd1 vccd1 _3447_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_2_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2653__A0 _2355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2500__S0 _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2239__A3 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3270_ _3484_/CLK _3270_/D vssd1 vssd1 vccd1 vccd1 _3270_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _2677_/B _2221_/B vssd1 vssd1 vccd1 vccd1 _2242_/C sky130_fd_sc_hd__or2_1
X_2152_ _2152_/A _2152_/B vssd1 vssd1 vccd1 vccd1 _2152_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__1686__A1 _2399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2083_ _3542_/Q _2084_/B vssd1 vssd1 vccd1 vccd1 _2083_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__2635__A0 _2358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2985_ _3110_/A vssd1 vssd1 vccd1 vccd1 _2985_/Y sky130_fd_sc_hd__inv_2
X_1936_ _1933_/Y _1934_/X _1935_/Y _1935_/B _1932_/A vssd1 vssd1 vccd1 vccd1 _1936_/X
+ sky130_fd_sc_hd__a32o_1
X_1867_ _1848_/A _1848_/B _1837_/A vssd1 vssd1 vccd1 vccd1 _1867_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout110_A hold126/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold811 _3545_/Q vssd1 vssd1 vccd1 vccd1 hold811/X sky130_fd_sc_hd__dlygate4sd3_1
X_1798_ _1791_/A _3150_/Q _1798_/C _1798_/D vssd1 vssd1 vccd1 vccd1 _1798_/X sky130_fd_sc_hd__and4b_1
X_3606_ _3607_/CLK _3606_/D _3097_/Y vssd1 vssd1 vccd1 vccd1 _3606_/Q sky130_fd_sc_hd__dfrtp_1
Xhold800 _3585_/Q vssd1 vssd1 vccd1 vccd1 hold800/X sky130_fd_sc_hd__dlygate4sd3_1
X_3537_ _3632_/CLK _3537_/D _3031_/Y vssd1 vssd1 vccd1 vccd1 _3537_/Q sky130_fd_sc_hd__dfrtp_1
Xhold855 _2332_/X vssd1 vssd1 vccd1 vccd1 _3383_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold844 _3542_/Q vssd1 vssd1 vccd1 vccd1 hold844/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold822 hold822/A vssd1 vssd1 vccd1 vccd1 _1941_/S sky130_fd_sc_hd__buf_1
Xhold833 _3550_/Q vssd1 vssd1 vccd1 vccd1 _1772_/B sky130_fd_sc_hd__buf_1
Xhold877 _2330_/X vssd1 vssd1 vccd1 vccd1 _3439_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 _3352_/Q vssd1 vssd1 vccd1 vccd1 _2144_/D sky130_fd_sc_hd__buf_1
Xhold888 _2198_/B vssd1 vssd1 vccd1 vccd1 _2375_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3468_ _3574_/CLK _3468_/D _2962_/Y vssd1 vssd1 vccd1 vccd1 _3468_/Q sky130_fd_sc_hd__dfrtp_1
Xhold899 _2257_/X vssd1 vssd1 vccd1 vccd1 _3464_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3399_ _3408_/CLK _3399_/D vssd1 vssd1 vccd1 vccd1 _3399_/Q sky130_fd_sc_hd__dfxtp_1
X_2419_ _3479_/Q _2507_/B _2417_/Y _2415_/X vssd1 vssd1 vccd1 vccd1 _2419_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2874__A0 _2109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2626__A0 _2098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2617__A0 _2109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2562__B hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2770_ _2800_/A _2790_/B vssd1 vssd1 vccd1 vccd1 _2779_/S sky130_fd_sc_hd__nor2_4
X_1721_ hold89/X _1845_/A vssd1 vssd1 vccd1 vccd1 _1721_/X sky130_fd_sc_hd__and2b_1
XANTENNA__1609__D input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1652_ _1569_/A _2400_/A hold53/X vssd1 vssd1 vccd1 vccd1 _3613_/D sky130_fd_sc_hd__mux2_1
Xhold107 _2418_/B vssd1 vssd1 vccd1 vccd1 _2413_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 _3308_/Q vssd1 vssd1 vccd1 vccd1 hold129/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 _1669_/X vssd1 vssd1 vccd1 vccd1 _3606_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1583_ _1847_/A vssd1 vssd1 vccd1 vccd1 _1583_/Y sky130_fd_sc_hd__inv_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _3322_/CLK _3322_/D vssd1 vssd1 vccd1 vccd1 _3322_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _3330_/CLK _3253_/D vssd1 vssd1 vccd1 vccd1 _3253_/Q sky130_fd_sc_hd__dfxtp_1
X_2204_ _2204_/A _2204_/B vssd1 vssd1 vccd1 vccd1 _2213_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_47_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3431_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3184_ _3433_/CLK _3184_/D vssd1 vssd1 vccd1 vccd1 _3184_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2856__A0 _2104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2135_ _2126_/A _2144_/C _2135_/C _2139_/B vssd1 vssd1 vccd1 vccd1 _2135_/X sky130_fd_sc_hd__and4b_1
XFILLER_0_88_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2608__A0 _2103_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2066_ _2096_/A _2084_/B vssd1 vssd1 vccd1 vccd1 _2067_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_76_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2968_ _3061_/A vssd1 vssd1 vccd1 vccd1 _2968_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2899__S _2900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1919_ _1912_/B _1918_/B _1935_/A vssd1 vssd1 vccd1 vccd1 _1919_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2899_ hold526/X _2073_/X _2900_/S vssd1 vssd1 vccd1 vccd1 _2899_/X sky130_fd_sc_hd__mux2_1
Xhold630 _3178_/Q vssd1 vssd1 vccd1 vccd1 hold630/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 _3392_/Q vssd1 vssd1 vccd1 vccd1 hold652/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 _2622_/X vssd1 vssd1 vccd1 vccd1 _3170_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold641 _2842_/X vssd1 vssd1 vccd1 vccd1 _3372_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 _3341_/Q vssd1 vssd1 vccd1 vccd1 hold674/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 _2874_/X vssd1 vssd1 vccd1 vccd1 _3405_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 _3371_/Q vssd1 vssd1 vccd1 vccd1 hold696/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2847__A0 _2357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1978__S _2000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1984__S1 _2219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2838__A0 _2355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2557__B hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2822_ hold510/X _2098_/S _2829_/S vssd1 vssd1 vccd1 vccd1 _2822_/X sky130_fd_sc_hd__mux2_1
X_2753_ hold339/X _2803_/A1 _2759_/S vssd1 vssd1 vccd1 vccd1 _2753_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1704_ _1704_/A _1704_/B vssd1 vssd1 vccd1 vccd1 _1704_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_41_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2684_ _2806_/A1 hold305/X _2687_/S vssd1 vssd1 vccd1 vccd1 _2684_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_53_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1635_ _3627_/Q hold45/X hold12/X vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__mux2_1
X_1566_ _2121_/A vssd1 vssd1 vccd1 vccd1 _2091_/S sky130_fd_sc_hd__inv_2
X_3305_ _3324_/CLK _3305_/D vssd1 vssd1 vccd1 vccd1 _3305_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _3326_/CLK _3236_/D vssd1 vssd1 vccd1 vccd1 _3236_/Q sky130_fd_sc_hd__dfxtp_1
X_3167_ _3433_/CLK _3167_/D vssd1 vssd1 vccd1 vccd1 _3167_/Q sky130_fd_sc_hd__dfxtp_1
X_3098_ _3112_/A vssd1 vssd1 vccd1 vccd1 _3098_/Y sky130_fd_sc_hd__inv_2
X_2118_ _1588_/Y _2117_/X _1811_/S vssd1 vssd1 vccd1 vccd1 _2118_/Y sky130_fd_sc_hd__a21oi_1
X_2049_ _3244_/Q _3316_/Q _3307_/Q _3298_/Q _2049_/S0 _2195_/A1 vssd1 vssd1 vccd1
+ vccd1 _2049_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_64_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout79 _1777_/C vssd1 vssd1 vccd1 vccd1 _2070_/A sky130_fd_sc_hd__clkbuf_8
Xfanout68 _1743_/Y vssd1 vssd1 vccd1 vccd1 _2387_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold471 _1911_/B vssd1 vssd1 vccd1 vccd1 hold471/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold460 _2226_/X vssd1 vssd1 vccd1 vccd1 _2227_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 _2817_/X vssd1 vssd1 vccd1 vccd1 _3340_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 _3584_/Q vssd1 vssd1 vccd1 vccd1 _2343_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2296__A1 hold59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3021_ _3032_/A vssd1 vssd1 vccd1 vccd1 _3021_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2805_ hold443/X _2805_/A1 _2809_/S vssd1 vssd1 vccd1 vccd1 _2805_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2736_ hold271/X _2806_/A1 _2739_/S vssd1 vssd1 vccd1 vccd1 _2736_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2667_ _2790_/A _2800_/B vssd1 vssd1 vccd1 vccd1 _2676_/S sky130_fd_sc_hd__nor2_4
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1618_ _1767_/S hold75/X _1622_/S vssd1 vssd1 vccd1 vccd1 _1618_/X sky130_fd_sc_hd__mux2_1
X_2598_ _2360_/B hold574/X _2601_/S vssd1 vssd1 vccd1 vccd1 _2598_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2197__B _2198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3219_ _3504_/CLK _3219_/D vssd1 vssd1 vccd1 vccd1 _3219_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3102__A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold290 _3199_/Q vssd1 vssd1 vccd1 vccd1 hold290/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3570_ _3571_/CLK _3570_/D _3064_/Y vssd1 vssd1 vccd1 vccd1 _3570_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2521_ _2520_/X _2517_/X _3518_/Q vssd1 vssd1 vccd1 vccd1 _2521_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2452_ _2451_/X _2448_/X _3518_/Q vssd1 vssd1 vccd1 vccd1 _2452_/X sky130_fd_sc_hd__mux2_1
X_2383_ _2383_/A _2383_/B vssd1 vssd1 vccd1 vccd1 _2911_/C sky130_fd_sc_hd__or2_1
XANTENNA_hold11_A hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput3 input3/A vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_2
X_3004_ _3110_/A vssd1 vssd1 vccd1 vccd1 _3004_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_74_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2719_ _2719_/A _2760_/A vssd1 vssd1 vccd1 vccd1 _2728_/S sky130_fd_sc_hd__or2_4
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2700__S _2707_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2671__A1 _2804_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2610__S _2612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2034__S0 _2045_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1952_ _2130_/B _2129_/A _2157_/A vssd1 vssd1 vccd1 vccd1 _2152_/A sky130_fd_sc_hd__and3_1
XFILLER_0_71_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1883_ _1883_/A _3523_/Q vssd1 vssd1 vccd1 vccd1 _1883_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3622_ _3622_/CLK _3622_/D _3113_/Y vssd1 vssd1 vccd1 vccd1 _3622_/Q sky130_fd_sc_hd__dfrtp_4
X_3553_ _3571_/CLK _3553_/D _3047_/Y vssd1 vssd1 vccd1 vccd1 _3553_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3484_ _3484_/CLK _3484_/D _2978_/Y vssd1 vssd1 vccd1 vccd1 _3484_/Q sky130_fd_sc_hd__dfrtp_1
X_2504_ _2503_/X _2502_/X _3517_/Q vssd1 vssd1 vccd1 vccd1 _2504_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2520__S _3517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2435_ _2435_/A _2575_/C vssd1 vssd1 vccd1 vccd1 _2508_/A sky130_fd_sc_hd__nor2_1
X_2366_ _1568_/Y _2105_/A _2365_/X vssd1 vssd1 vccd1 vccd1 _2367_/C sky130_fd_sc_hd__o21ba_1
X_2297_ _1730_/B _2406_/A hold22/X vssd1 vssd1 vccd1 vccd1 _3448_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_78_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2500__S1 _1943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2016__S0 _2221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2605__S _2612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _2677_/B _2221_/B vssd1 vssd1 vccd1 vccd1 _2242_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_17_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2576__A _2576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2151_ _1955_/D _2133_/C _2158_/S _2150_/X _2130_/A vssd1 vssd1 vccd1 vccd1 _2151_/Y
+ sky130_fd_sc_hd__o32ai_1
X_2082_ _2092_/A _2080_/Y _2081_/Y vssd1 vssd1 vccd1 vccd1 _2082_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_88_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2984_ _3097_/A vssd1 vssd1 vccd1 vccd1 _2984_/Y sky130_fd_sc_hd__inv_2
X_1935_ _1935_/A _1935_/B vssd1 vssd1 vccd1 vccd1 _1935_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_83_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2494__S0 _2532_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1866_ _1837_/A _1849_/Y _1865_/X _1865_/A _1836_/A vssd1 vssd1 vccd1 vccd1 _1866_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_71_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3605_ _3605_/CLK _3605_/D _3096_/Y vssd1 vssd1 vccd1 vccd1 _3605_/Q sky130_fd_sc_hd__dfrtp_1
Xhold812 _1830_/X vssd1 vssd1 vccd1 vccd1 _3544_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1797_ _1600_/Y _1798_/C _1798_/D vssd1 vssd1 vccd1 vccd1 _1801_/A sky130_fd_sc_hd__o21ai_1
Xhold801 _2368_/X vssd1 vssd1 vccd1 vccd1 _3343_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3536_ _3632_/CLK _3536_/D _3030_/Y vssd1 vssd1 vccd1 vccd1 _3536_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold823 _3470_/Q vssd1 vssd1 vccd1 vccd1 _2248_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold845 _1832_/X vssd1 vssd1 vccd1 vccd1 _3542_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout103_A hold87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2020__C1 _2000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold834 _1805_/Y vssd1 vssd1 vccd1 vccd1 hold834/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 _2227_/A vssd1 vssd1 vccd1 vccd1 _2193_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 _3464_/Q vssd1 vssd1 vccd1 vccd1 hold878/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 _3514_/Q vssd1 vssd1 vccd1 vccd1 _1932_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold867 _2378_/X vssd1 vssd1 vccd1 vccd1 _3352_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3467_ _3575_/CLK _3467_/D _2961_/Y vssd1 vssd1 vccd1 vccd1 _3467_/Q sky130_fd_sc_hd__dfrtp_1
X_3398_ _3434_/CLK _3398_/D vssd1 vssd1 vccd1 vccd1 _3398_/Q sky130_fd_sc_hd__dfxtp_1
X_2418_ hold9/A _2418_/B vssd1 vssd1 vccd1 vccd1 _2507_/B sky130_fd_sc_hd__or2_2
X_2349_ _2349_/A _2349_/B vssd1 vssd1 vccd1 vccd1 _2349_/X sky130_fd_sc_hd__or2_1
XFILLER_0_79_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2865__A1 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xuart_macro_wrapper_130 vssd1 vssd1 vccd1 vccd1 uart_macro_wrapper_130/HI io_oeb[1]
+ sky130_fd_sc_hd__conb_1
X_1720_ _1871_/A hold73/X vssd1 vssd1 vccd1 vccd1 _1720_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1651_ _1568_/A _2401_/A hold53/X vssd1 vssd1 vccd1 vccd1 _3614_/D sky130_fd_sc_hd__mux2_1
Xhold108 _2437_/B vssd1 vssd1 vccd1 vccd1 _2576_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold119 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 input28/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1582_ _1850_/A vssd1 vssd1 vccd1 vccd1 _1582_/Y sky130_fd_sc_hd__inv_2
X_3321_ _3321_/CLK _3321_/D vssd1 vssd1 vccd1 vccd1 _3321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _3324_/CLK _3252_/D vssd1 vssd1 vccd1 vccd1 _3252_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2203_ _3479_/Q _2215_/B vssd1 vssd1 vccd1 vccd1 _2204_/B sky130_fd_sc_hd__nand2_1
X_3183_ _3434_/CLK _3183_/D vssd1 vssd1 vccd1 vccd1 _3183_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2134_ _2000_/S _2135_/C _2139_/B vssd1 vssd1 vccd1 vccd1 _2138_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2065_ _2065_/A _2065_/B vssd1 vssd1 vccd1 vccd1 _2065_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_16_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3605_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2967_ _3061_/A vssd1 vssd1 vccd1 vccd1 _2967_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2467__S0 _2532_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2898_ hold498/X _2072_/Y _2900_/S vssd1 vssd1 vccd1 vccd1 _2898_/X sky130_fd_sc_hd__mux2_1
X_1918_ _1911_/B _1918_/B vssd1 vssd1 vccd1 vccd1 _1918_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_32_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1849_ _1865_/A _1865_/B vssd1 vssd1 vccd1 vccd1 _1849_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold620 _3166_/Q vssd1 vssd1 vccd1 vccd1 hold620/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 _2859_/X vssd1 vssd1 vccd1 vccd1 _3392_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold642 _3424_/Q vssd1 vssd1 vccd1 vccd1 hold642/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 _2631_/X vssd1 vssd1 vccd1 vccd1 _3178_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 _2818_/X vssd1 vssd1 vccd1 vccd1 _3341_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 _2841_/X vssd1 vssd1 vccd1 vccd1 _3371_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 _3406_/Q vssd1 vssd1 vccd1 vccd1 hold664/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 _3194_/Q vssd1 vssd1 vccd1 vccd1 hold686/X sky130_fd_sc_hd__dlygate4sd3_1
X_3519_ _3521_/CLK _3519_/D _3013_/Y vssd1 vssd1 vccd1 vccd1 _3519_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2783__A0 _2803_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2821_ hold528/X _2358_/B _2829_/S vssd1 vssd1 vccd1 vccd1 _2821_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2449__S0 _2532_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2752_ hold140/X _2802_/A1 _2759_/S vssd1 vssd1 vccd1 vccd1 _2752_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1703_ _1700_/B hold885/X _3462_/D vssd1 vssd1 vccd1 vccd1 _1703_/Y sky130_fd_sc_hd__a21oi_1
X_2683_ _2805_/A1 hold431/X _2687_/S vssd1 vssd1 vccd1 vccd1 _2683_/X sky130_fd_sc_hd__mux2_1
X_1634_ _1560_/A _2406_/A hold12/X vssd1 vssd1 vccd1 vccd1 _3628_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1565_ _2070_/A vssd1 vssd1 vccd1 vccd1 _2058_/C sky130_fd_sc_hd__inv_2
X_3304_ _3322_/CLK _3304_/D vssd1 vssd1 vccd1 vccd1 _3304_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3235_ _3329_/CLK _3235_/D vssd1 vssd1 vccd1 vccd1 _3235_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2829__A1 _2356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3166_ _3433_/CLK _3166_/D vssd1 vssd1 vccd1 vccd1 _3166_/Q sky130_fd_sc_hd__dfxtp_1
X_2117_ _2112_/X _2113_/X _2116_/X _1769_/B _1601_/Y vssd1 vssd1 vccd1 vccd1 _2117_/X
+ sky130_fd_sc_hd__a311o_1
X_3097_ _3097_/A vssd1 vssd1 vccd1 vccd1 _3097_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_55_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2048_ _3289_/Q _3280_/Q _3271_/Q _3262_/Q _2049_/S0 _2219_/A vssd1 vssd1 vccd1 vccd1
+ _2048_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2462__C1 _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout69 _2108_/Y vssd1 vssd1 vccd1 vccd1 _2109_/B sky130_fd_sc_hd__buf_4
XANTENNA__2703__S _2707_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2765__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold472 _1949_/X vssd1 vssd1 vccd1 vccd1 _3510_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold450 _2672_/X vssd1 vssd1 vccd1 vccd1 _3212_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 _2227_/X vssd1 vssd1 vccd1 vccd1 _3478_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _3402_/Q vssd1 vssd1 vccd1 vccd1 hold494/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 _2343_/Y vssd1 vssd1 vccd1 vccd1 _3346_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout83_A _2532_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1989__S _2000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3020_ _3061_/A vssd1 vssd1 vccd1 vccd1 _3020_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_73_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2804_ hold243/X _2804_/A1 _2809_/S vssd1 vssd1 vccd1 vccd1 _2804_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2747__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2735_ hold276/X _2805_/A1 _2739_/S vssd1 vssd1 vccd1 vccd1 _2735_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2666_ _2406_/A hold399/X _2666_/S vssd1 vssd1 vccd1 vccd1 _2666_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1617_ _2289_/A _2572_/A vssd1 vssd1 vccd1 vccd1 _1622_/S sky130_fd_sc_hd__nor2_2
X_2597_ _2104_/B hold568/X _2601_/S vssd1 vssd1 vccd1 vccd1 _2597_/X sky130_fd_sc_hd__mux2_1
X_3218_ _3333_/CLK _3218_/D vssd1 vssd1 vccd1 vccd1 _3218_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_31_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3627_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3149_ _3550_/CLK _3149_/D _2913_/Y vssd1 vssd1 vccd1 vccd1 _3149_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2433__S _3518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold280 _3321_/Q vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2910__A0 _2356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold291 _2658_/X vssd1 vssd1 vccd1 vccd1 _3199_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2608__S _2612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2426__C1 _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2520_ _2519_/X _2518_/X _3517_/Q vssd1 vssd1 vccd1 vccd1 _2520_/X sky130_fd_sc_hd__mux2_1
X_2451_ _2450_/X _2449_/X _2546_/S vssd1 vssd1 vccd1 vccd1 _2451_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2382_ _2000_/S _2377_/X hold986/X _1599_/Y vssd1 vssd1 vccd1 vccd1 _2382_/Y sky130_fd_sc_hd__o22ai_1
Xinput4 input4/A vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_2
X_3003_ _3110_/A vssd1 vssd1 vccd1 vccd1 _3003_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1658__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2718_ _2406_/A hold357/X _2718_/S vssd1 vssd1 vccd1 vccd1 _2718_/X sky130_fd_sc_hd__mux2_1
X_2649_ _2105_/A hold730/X _2654_/S vssd1 vssd1 vccd1 vccd1 _2649_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2952__A _3124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2399__A _2399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2034__S1 _2045_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1951_ _2129_/A _3492_/Q vssd1 vssd1 vccd1 vccd1 _2155_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1882_ _1837_/A _1879_/B _1881_/X _1839_/A _1836_/A vssd1 vssd1 vccd1 vccd1 _1882_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3621_ _3622_/CLK _3621_/D _3112_/Y vssd1 vssd1 vccd1 vccd1 _3621_/Q sky130_fd_sc_hd__dfrtp_1
X_3552_ _3571_/CLK _3552_/D _3046_/Y vssd1 vssd1 vccd1 vccd1 _3552_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2503_ _3177_/Q _3426_/Q _3417_/Q _3159_/Q _1918_/B _2532_/S1 vssd1 vssd1 vccd1 vccd1
+ _2503_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3483_ _3605_/CLK _3483_/D _2977_/Y vssd1 vssd1 vccd1 vccd1 _3483_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2434_ _1908_/D _2433_/X _2426_/X vssd1 vssd1 vccd1 vccd1 _2434_/X sky130_fd_sc_hd__a21o_2
X_2365_ _1568_/Y _2105_/A _2103_/Y _1567_/Y vssd1 vssd1 vccd1 vccd1 _2365_/X sky130_fd_sc_hd__a22o_1
X_2296_ _3449_/Q hold59/X hold22/X vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__mux2_1
XFILLER_0_78_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2711__S _2718_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3108__A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2016__S1 _2219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2150_ _2152_/A _2157_/B _2148_/B _2375_/A vssd1 vssd1 vccd1 vccd1 _2150_/X sky130_fd_sc_hd__o211a_1
X_2081_ _2092_/A _3540_/Q _2065_/A vssd1 vssd1 vccd1 vccd1 _2081_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2983_ _3097_/A vssd1 vssd1 vccd1 vccd1 _2983_/Y sky130_fd_sc_hd__inv_2
X_1934_ _1934_/A _1934_/B _1934_/C vssd1 vssd1 vccd1 vccd1 _1934_/X sky130_fd_sc_hd__or3_1
XFILLER_0_83_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2494__S1 _2532_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1865_ _1865_/A _1865_/B vssd1 vssd1 vccd1 vccd1 _1865_/X sky130_fd_sc_hd__or2_1
XFILLER_0_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold802 _3546_/Q vssd1 vssd1 vccd1 vccd1 hold802/X sky130_fd_sc_hd__dlygate4sd3_1
X_1796_ _1600_/Y _2387_/C _1795_/Y _2383_/A _3150_/D vssd1 vssd1 vccd1 vccd1 _1798_/D
+ sky130_fd_sc_hd__o221a_2
X_3604_ _3607_/CLK _3604_/D _3095_/Y vssd1 vssd1 vccd1 vccd1 _3604_/Q sky130_fd_sc_hd__dfrtp_1
X_3535_ _3632_/CLK _3535_/D _3029_/Y vssd1 vssd1 vccd1 vccd1 _3535_/Q sky130_fd_sc_hd__dfrtp_1
Xhold824 _2251_/X vssd1 vssd1 vccd1 vccd1 _3470_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 _3471_/Q vssd1 vssd1 vccd1 vccd1 hold846/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold813 _3539_/Q vssd1 vssd1 vccd1 vccd1 hold813/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 _1806_/Y vssd1 vssd1 vccd1 vccd1 _3552_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold868 _3474_/Q vssd1 vssd1 vccd1 vccd1 _2259_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 _2256_/X vssd1 vssd1 vccd1 vccd1 _3465_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3466_ _3575_/CLK _3466_/D _2960_/Y vssd1 vssd1 vccd1 vccd1 _3466_/Q sky130_fd_sc_hd__dfrtp_1
Xhold857 _1936_/X vssd1 vssd1 vccd1 vccd1 _3514_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2417_ _1924_/A _2575_/C _2435_/A vssd1 vssd1 vccd1 vccd1 _2417_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3397_ _3433_/CLK _3397_/D vssd1 vssd1 vccd1 vccd1 _3397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2348_ _1596_/Y _2347_/X hold478/X vssd1 vssd1 vccd1 vccd1 _2348_/Y sky130_fd_sc_hd__a21oi_1
X_2279_ _2271_/B _2281_/B _2283_/A vssd1 vssd1 vccd1 vccd1 _2279_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2706__S _2707_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xuart_macro_wrapper_131 vssd1 vssd1 vccd1 vccd1 uart_macro_wrapper_131/HI wbs_dat_o[17]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_80_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1650_ _3615_/Q hold75/X hold53/X vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__mux2_1
X_1581_ _1851_/A vssd1 vssd1 vccd1 vccd1 _1581_/Y sky130_fd_sc_hd__inv_2
Xhold109 _2576_/X vssd1 vssd1 vccd1 vccd1 _3591_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3320_ _3320_/CLK _3320_/D vssd1 vssd1 vccd1 vccd1 _3320_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2305__A1 _2576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3251_ _3324_/CLK _3251_/D vssd1 vssd1 vccd1 vccd1 _3251_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2202_ _2202_/A _2208_/B vssd1 vssd1 vccd1 vccd1 _2215_/B sky130_fd_sc_hd__xnor2_1
X_3182_ _3431_/CLK _3182_/D vssd1 vssd1 vccd1 vccd1 _3182_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2133_ _2379_/B _2133_/B _2133_/C _2133_/D vssd1 vssd1 vccd1 vccd1 _2139_/B sky130_fd_sc_hd__and4_2
X_2064_ _2064_/A _2064_/B vssd1 vssd1 vccd1 vccd1 _2090_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_44_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2966_ _3097_/A vssd1 vssd1 vccd1 vccd1 _2966_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2467__S1 _1912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2897_ hold512/X _2106_/X _2900_/S vssd1 vssd1 vccd1 vccd1 _2897_/X sky130_fd_sc_hd__mux2_1
X_1917_ _2546_/S hold471/X _1911_/Y _2160_/B vssd1 vssd1 vccd1 vccd1 _3517_/D sky130_fd_sc_hd__a22o_1
X_1848_ _1848_/A _1848_/B vssd1 vssd1 vccd1 vccd1 _1865_/B sky130_fd_sc_hd__and2_1
XANTENNA__2792__A1 _2802_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold610 _3357_/Q vssd1 vssd1 vccd1 vccd1 hold610/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold621 _2618_/X vssd1 vssd1 vccd1 vccd1 _3166_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold632 _3387_/Q vssd1 vssd1 vccd1 vccd1 hold632/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 _3434_/Q vssd1 vssd1 vccd1 vccd1 hold654/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold643 _2895_/X vssd1 vssd1 vccd1 vccd1 _3424_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1779_ _2092_/A _2096_/A vssd1 vssd1 vccd1 vccd1 _2123_/A sky130_fd_sc_hd__or2_1
Xhold676 _3420_/Q vssd1 vssd1 vccd1 vccd1 hold676/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 _2875_/X vssd1 vssd1 vccd1 vccd1 _3406_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 _2650_/X vssd1 vssd1 vccd1 vccd1 _3194_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3518_ _3614_/CLK _3518_/D _3012_/Y vssd1 vssd1 vccd1 vccd1 _3518_/Q sky130_fd_sc_hd__dfrtp_4
X_3449_ _3589_/CLK hold60/X _2943_/Y vssd1 vssd1 vccd1 vccd1 _3449_/Q sky130_fd_sc_hd__dfrtp_1
Xhold698 _3140_/Q vssd1 vssd1 vccd1 vccd1 hold698/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3121__A _3124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1969__S0 _2045_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2046__A_N _2036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2449__S1 _2532_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2820_ _2891_/A _2830_/B vssd1 vssd1 vccd1 vccd1 _2829_/S sky130_fd_sc_hd__and2_4
XFILLER_0_38_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2751_ hold245/X _2801_/A1 _2759_/S vssd1 vssd1 vccd1 vccd1 _2751_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1702_ _1702_/A _1702_/B vssd1 vssd1 vccd1 vccd1 _1702_/Y sky130_fd_sc_hd__nand2_1
X_2682_ _2804_/A1 hold237/X _2687_/S vssd1 vssd1 vccd1 vccd1 _2682_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_53_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2774__A1 _2804_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1633_ hold67/X hold59/X hold12/X vssd1 vssd1 vccd1 vccd1 _3629_/D sky130_fd_sc_hd__mux2_1
X_1564_ _3623_/Q vssd1 vssd1 vccd1 vccd1 _1564_/Y sky130_fd_sc_hd__inv_2
X_3303_ _3321_/CLK _3303_/D vssd1 vssd1 vccd1 vccd1 _3303_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _3408_/CLK _3234_/D vssd1 vssd1 vccd1 vccd1 _3234_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3165_ _3434_/CLK _3165_/D vssd1 vssd1 vccd1 vccd1 _3165_/Q sky130_fd_sc_hd__dfxtp_1
X_3096_ _3124_/A vssd1 vssd1 vccd1 vccd1 _3096_/Y sky130_fd_sc_hd__inv_2
X_2116_ _2116_/A hold99/X _2116_/C _2116_/D vssd1 vssd1 vccd1 vccd1 _2116_/X sky130_fd_sc_hd__or4_1
X_2047_ _3217_/Q _3208_/Q _3199_/Q _3325_/Q _3483_/Q _2195_/A1 vssd1 vssd1 vccd1 vccd1
+ _2047_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_49_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2949_ _3122_/A vssd1 vssd1 vccd1 vccd1 _2949_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold451 _3622_/Q vssd1 vssd1 vccd1 vccd1 _2063_/A sky130_fd_sc_hd__clkbuf_2
Xhold440 _2663_/X vssd1 vssd1 vccd1 vccd1 _3204_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 _3488_/Q vssd1 vssd1 vccd1 vccd1 _2176_/A sky130_fd_sc_hd__buf_1
Xhold495 _2870_/X vssd1 vssd1 vccd1 vccd1 _3402_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 _3510_/Q vssd1 vssd1 vccd1 vccd1 _1923_/A sky130_fd_sc_hd__clkbuf_2
Xhold484 _3587_/Q vssd1 vssd1 vccd1 vccd1 _2336_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2453__B1 _2445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2756__A1 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_1_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3329_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_58_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2803_ hold382/X _2803_/A1 _2809_/S vssd1 vssd1 vccd1 vccd1 _2803_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2105__A _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2734_ hold167/X _2804_/A1 _2739_/S vssd1 vssd1 vccd1 vccd1 _2734_/X sky130_fd_sc_hd__mux2_1
X_2665_ _2808_/A1 hold212/X _2666_/S vssd1 vssd1 vccd1 vccd1 _2665_/X sky130_fd_sc_hd__mux2_1
X_2596_ _2105_/A hold562/X _2601_/S vssd1 vssd1 vccd1 vccd1 _2596_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1616_ hold35/X hold94/X vssd1 vssd1 vccd1 vccd1 _2572_/A sky130_fd_sc_hd__nand2_2
X_3217_ _3330_/CLK _3217_/D vssd1 vssd1 vccd1 vccd1 _3217_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2683__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3148_ _3576_/CLK _3148_/D _1605_/Y vssd1 vssd1 vccd1 vccd1 _3148_/Q sky130_fd_sc_hd__dfstp_1
X_3079_ _3090_/A vssd1 vssd1 vccd1 vccd1 _3079_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2714__S _2718_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2738__A1 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold270 _2771_/X vssd1 vssd1 vccd1 vccd1 _3298_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 _2796_/X vssd1 vssd1 vccd1 vccd1 _3321_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _3208_/Q vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2450_ _3173_/Q _3422_/Q _3413_/Q _3155_/Q _2532_/S0 _1912_/B vssd1 vssd1 vccd1 vccd1
+ _2450_/X sky130_fd_sc_hd__mux4_1
X_2381_ _2381_/A _2381_/B _2381_/C _2381_/D vssd1 vssd1 vccd1 vccd1 _2381_/X sky130_fd_sc_hd__or4_1
Xinput5 input5/A vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_1
X_3002_ _3110_/A vssd1 vssd1 vccd1 vccd1 _3002_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2665__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2534__S _3518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1640__A1 _2400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout126_A _3057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2717_ _2808_/A1 hold218/X _2718_/S vssd1 vssd1 vccd1 vccd1 _2717_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1674__A hold62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2648_ _2109_/B hold540/X _2654_/S vssd1 vssd1 vccd1 vccd1 _2648_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2579_ _2729_/B _2708_/A vssd1 vssd1 vccd1 vccd1 _2719_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_84_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2503__S0 _1918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1631__A1 hold78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2647__A0 _2098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1950_ _1950_/A _1950_/B _1950_/C vssd1 vssd1 vccd1 vccd1 _2379_/B sky130_fd_sc_hd__and3_1
X_1881_ _1883_/A _3523_/Q _1839_/A vssd1 vssd1 vccd1 vccd1 _1881_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_28_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1622__A1 _2576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3620_ _3627_/CLK _3620_/D _3111_/Y vssd1 vssd1 vccd1 vccd1 _3620_/Q sky130_fd_sc_hd__dfrtp_1
X_3551_ _3559_/CLK _3551_/D _3045_/Y vssd1 vssd1 vccd1 vccd1 _3551_/Q sky130_fd_sc_hd__dfrtp_1
X_2502_ _3376_/Q _3358_/Q _3367_/Q _3195_/Q _1918_/B _1912_/B vssd1 vssd1 vccd1 vccd1
+ _2502_/X sky130_fd_sc_hd__mux4_1
X_3482_ _3605_/CLK _3482_/D _2976_/Y vssd1 vssd1 vccd1 vccd1 _3482_/Q sky130_fd_sc_hd__dfrtp_1
X_2433_ _2432_/X _2429_/X _3518_/Q vssd1 vssd1 vccd1 vccd1 _2433_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2886__A0 _2104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2364_ _1570_/Y _2098_/S _2109_/B _1569_/Y _2363_/X vssd1 vssd1 vccd1 vccd1 _2367_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2295_ _3450_/Q hold5/X hold22/A vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__mux2_1
XANTENNA__2638__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2877__A0 _2360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3124__A _3124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2629__A0 _2103_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1745__C _1769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2080_ _3541_/Q _2084_/B vssd1 vssd1 vccd1 vccd1 _2080_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2982_ _3097_/A vssd1 vssd1 vccd1 vccd1 _2982_/Y sky130_fd_sc_hd__inv_2
X_1933_ _1934_/A _1934_/B _1934_/C vssd1 vssd1 vccd1 vccd1 _1933_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1864_ _1863_/X _1851_/B _1850_/A _1836_/A vssd1 vssd1 vccd1 vccd1 _3534_/D sky130_fd_sc_hd__a2bb2o_1
X_3603_ _3605_/CLK _3603_/D _3094_/Y vssd1 vssd1 vccd1 vccd1 _3603_/Q sky130_fd_sc_hd__dfrtp_1
Xinput30 hold74/X vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__buf_1
XFILLER_0_12_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold803 _1829_/X vssd1 vssd1 vccd1 vccd1 _3545_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1795_ _1809_/A _1795_/B vssd1 vssd1 vccd1 vccd1 _1795_/Y sky130_fd_sc_hd__nand2_1
X_3534_ _3632_/CLK _3534_/D _3028_/Y vssd1 vssd1 vccd1 vccd1 _3534_/Q sky130_fd_sc_hd__dfrtp_1
Xhold825 _3475_/Q vssd1 vssd1 vccd1 vccd1 _2259_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 _1835_/X vssd1 vssd1 vccd1 vccd1 _3539_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold836 _3547_/Q vssd1 vssd1 vccd1 vccd1 hold836/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 _2237_/Y vssd1 vssd1 vccd1 vccd1 _2238_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3465_ _3574_/CLK _3465_/D _2959_/Y vssd1 vssd1 vccd1 vccd1 _3465_/Q sky130_fd_sc_hd__dfrtp_1
Xhold858 _3468_/Q vssd1 vssd1 vccd1 vccd1 hold858/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 _2250_/X vssd1 vssd1 vccd1 vccd1 _3471_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2859__A0 _2355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2416_ _2416_/A hold20/X vssd1 vssd1 vccd1 vccd1 _2575_/C sky130_fd_sc_hd__and2_1
X_3396_ _3432_/CLK _3396_/D vssd1 vssd1 vccd1 vccd1 _3396_/Q sky130_fd_sc_hd__dfxtp_1
X_2347_ _1575_/Y _2208_/A _2345_/X _2346_/X hold459/X vssd1 vssd1 vccd1 vccd1 _2347_/X
+ sky130_fd_sc_hd__a221o_1
X_2278_ _2283_/A _2278_/B _2278_/C vssd1 vssd1 vccd1 vccd1 _2278_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__2722__S _2728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2011__A1 _2144_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2632__S _2633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuart_macro_wrapper_132 vssd1 vssd1 vccd1 vccd1 uart_macro_wrapper_132/HI wbs_dat_o[20]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_80_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1580_ _1855_/A vssd1 vssd1 vccd1 vccd1 _1580_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2553__A2 hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3590_/CLK _3250_/D vssd1 vssd1 vccd1 vccd1 _3250_/Q sky130_fd_sc_hd__dfxtp_1
X_2201_ _2202_/A _2205_/B vssd1 vssd1 vccd1 vccd1 _2204_/A sky130_fd_sc_hd__nand2_1
X_3181_ _3432_/CLK _3181_/D vssd1 vssd1 vccd1 vccd1 _3181_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2132_ _2146_/A _2379_/C _2144_/C vssd1 vssd1 vccd1 vccd1 _2133_/D sky130_fd_sc_hd__mux2_1
X_2063_ _2063_/A _2070_/A vssd1 vssd1 vccd1 vccd1 _2065_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_88_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2965_ _3069_/A vssd1 vssd1 vccd1 vccd1 _2965_/Y sky130_fd_sc_hd__inv_2
X_2896_ hold542/X _2104_/B _2900_/S vssd1 vssd1 vccd1 vccd1 _2896_/X sky130_fd_sc_hd__mux2_1
X_1916_ _1916_/A _1916_/B vssd1 vssd1 vccd1 vccd1 _2160_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1847_ _1847_/A _1871_/A _1871_/B vssd1 vssd1 vccd1 vccd1 _1848_/B sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_25_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3567_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold600 _3365_/Q vssd1 vssd1 vccd1 vccd1 hold600/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 _2825_/X vssd1 vssd1 vccd1 vccd1 _3357_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 _3364_/Q vssd1 vssd1 vccd1 vccd1 hold644/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 _2854_/X vssd1 vssd1 vccd1 vccd1 _3387_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold622 _3173_/Q vssd1 vssd1 vccd1 vccd1 hold622/X sky130_fd_sc_hd__dlygate4sd3_1
X_3517_ _3614_/CLK _3517_/D _3011_/Y vssd1 vssd1 vccd1 vccd1 _3517_/Q sky130_fd_sc_hd__dfrtp_4
X_1778_ _2121_/A _2096_/A vssd1 vssd1 vccd1 vccd1 _2319_/A sky130_fd_sc_hd__nor2_1
Xhold655 _2906_/X vssd1 vssd1 vccd1 vccd1 _3434_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 _2890_/X vssd1 vssd1 vccd1 vccd1 _3420_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 _3410_/Q vssd1 vssd1 vccd1 vccd1 hold688/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 _3187_/Q vssd1 vssd1 vccd1 vccd1 hold666/X sky130_fd_sc_hd__dlygate4sd3_1
X_3448_ _3633_/CLK _3448_/D _2942_/Y vssd1 vssd1 vccd1 vccd1 _3448_/Q sky130_fd_sc_hd__dfrtp_1
Xhold699 _2594_/X vssd1 vssd1 vccd1 vccd1 _3140_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ _3516_/CLK _3379_/D vssd1 vssd1 vccd1 vccd1 _3379_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2717__S _2718_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_3__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2452__S _3518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__1969__S1 _2045_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2299__A1 hold87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2627__S _2633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2750_ _2790_/A _2760_/B vssd1 vssd1 vccd1 vccd1 _2759_/S sky130_fd_sc_hd__nor2_4
XFILLER_0_5_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1701_ _1698_/B hold893/X _3462_/D vssd1 vssd1 vccd1 vccd1 _1701_/Y sky130_fd_sc_hd__a21oi_1
X_2681_ _2803_/A1 hold378/X _2687_/S vssd1 vssd1 vccd1 vccd1 _2681_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1632_ _3630_/Q hold5/X hold12/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1563_ _2387_/A vssd1 vssd1 vccd1 vccd1 _2490_/A sky130_fd_sc_hd__inv_2
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3302_ _3320_/CLK _3302_/D vssd1 vssd1 vccd1 vccd1 _3302_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _3332_/CLK _3233_/D vssd1 vssd1 vccd1 vccd1 _3233_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3164_ _3434_/CLK _3164_/D vssd1 vssd1 vccd1 vccd1 _3164_/Q sky130_fd_sc_hd__dfxtp_1
X_2115_ hold72/X _2383_/B vssd1 vssd1 vccd1 vccd1 _2116_/D sky130_fd_sc_hd__nor2_1
X_3095_ _3097_/A vssd1 vssd1 vccd1 vccd1 _3095_/Y sky130_fd_sc_hd__inv_2
X_2046_ _2036_/S _2046_/B vssd1 vssd1 vccd1 vccd1 _2046_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_71_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2948_ _3122_/A vssd1 vssd1 vccd1 vccd1 _2948_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2879_ _2355_/B hold688/X _2880_/S vssd1 vssd1 vccd1 vccd1 _2879_/X sky130_fd_sc_hd__mux2_1
Xhold452 _3628_/Q vssd1 vssd1 vccd1 vccd1 _1560_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 _3479_/Q vssd1 vssd1 vccd1 vccd1 _2217_/S sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold430 _2674_/X vssd1 vssd1 vccd1 vccd1 _3214_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 _3203_/Q vssd1 vssd1 vccd1 vccd1 hold441/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 _3356_/Q vssd1 vssd1 vccd1 vccd1 hold496/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 _1932_/B vssd1 vssd1 vccd1 vccd1 _1929_/B sky130_fd_sc_hd__buf_1
Xhold485 _2336_/Y vssd1 vssd1 vccd1 vccd1 _3381_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2453__A1 _1908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1753__C _1769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2692__A1 _2804_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2802_ hold174/X _2802_/A1 _2809_/S vssd1 vssd1 vccd1 vccd1 _2802_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2733_ hold334/X _2803_/A1 _2739_/S vssd1 vssd1 vccd1 vccd1 _2733_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2664_ _2807_/A1 hold427/X _2666_/S vssd1 vssd1 vccd1 vccd1 _2664_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2595_ _2109_/B hold710/X _2601_/S vssd1 vssd1 vccd1 vccd1 _2595_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1944__B _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1615_ hold35/A hold94/A vssd1 vssd1 vccd1 vccd1 _2510_/A sky130_fd_sc_hd__and2_2
XFILLER_0_5_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3216_ _3333_/CLK _3216_/D vssd1 vssd1 vccd1 vccd1 _3216_/Q sky130_fd_sc_hd__dfxtp_1
X_3147_ _3432_/CLK _3147_/D vssd1 vssd1 vccd1 vccd1 _3147_/Q sky130_fd_sc_hd__dfxtp_1
X_3078_ _3090_/A vssd1 vssd1 vccd1 vccd1 _3078_/Y sky130_fd_sc_hd__inv_2
X_2029_ _2028_/X _2027_/X _2222_/A vssd1 vssd1 vccd1 vccd1 _2029_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_49_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_40_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3413_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold260 _2781_/X vssd1 vssd1 vccd1 vccd1 _3307_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 _3267_/Q vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _3285_/Q vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 _2668_/X vssd1 vssd1 vccd1 vccd1 _3208_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2674__A1 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2037__S0 _2221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2362__B1 _2109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2380_ _2144_/A _2372_/S hold904/X _2387_/A vssd1 vssd1 vccd1 vccd1 _2380_/X sky130_fd_sc_hd__a22o_1
Xinput6 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3001_ _3101_/A vssd1 vssd1 vccd1 vccd1 _3001_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1658__C input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2716_ _2807_/A1 hold359/X _2718_/S vssd1 vssd1 vccd1 vccd1 _2716_/X sky130_fd_sc_hd__mux2_1
X_2647_ _2098_/S hold734/X _2654_/S vssd1 vssd1 vccd1 vccd1 _2647_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout119_A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2578_ _3488_/Q _2578_/B vssd1 vssd1 vccd1 vccd1 _2790_/A sky130_fd_sc_hd__nand2b_4
XFILLER_0_77_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2725__S _2728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2503__S1 _2532_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2895__A1 _2101_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ _1837_/A _1841_/Y _1879_/Y _1840_/A _1836_/A vssd1 vssd1 vccd1 vccd1 _1880_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3550_ _3550_/CLK _3550_/D _3044_/Y vssd1 vssd1 vccd1 vccd1 _3550_/Q sky130_fd_sc_hd__dfrtp_1
X_2501_ _2500_/X _2499_/X _2546_/S vssd1 vssd1 vccd1 vccd1 _2501_/X sky130_fd_sc_hd__mux2_1
X_3481_ _3605_/CLK _3481_/D _2975_/Y vssd1 vssd1 vccd1 vccd1 _3481_/Q sky130_fd_sc_hd__dfrtp_1
X_2432_ _2431_/X _2430_/X _2546_/S vssd1 vssd1 vccd1 vccd1 _2432_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2430__S0 _1918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2363_ _2363_/A _2363_/B _2363_/C _2363_/D vssd1 vssd1 vccd1 vccd1 _2363_/X sky130_fd_sc_hd__and4_1
XFILLER_0_47_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2294_ _3451_/Q hold78/X hold22/X vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__mux2_1
XFILLER_0_2_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2497__S0 _3517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2801__A1 _2801_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2868__A1 _2357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1761__C _1769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2981_ _3097_/A vssd1 vssd1 vccd1 vccd1 _2981_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_56_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1932_ _1932_/A _1932_/B vssd1 vssd1 vccd1 vccd1 _1934_/C sky130_fd_sc_hd__xor2_1
X_1863_ _1582_/Y _1849_/Y _1837_/Y vssd1 vssd1 vccd1 vccd1 _1863_/X sky130_fd_sc_hd__a21o_1
Xinput20 input20/A vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_1
X_3602_ _3602_/CLK _3602_/D _3093_/Y vssd1 vssd1 vccd1 vccd1 _3602_/Q sky130_fd_sc_hd__dfrtp_1
Xinput31 hold69/X vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__buf_1
XFILLER_0_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1794_ _1809_/A _1773_/Y _1793_/Y _1825_/A vssd1 vssd1 vccd1 vccd1 _1794_/X sky130_fd_sc_hd__a22o_1
X_3533_ _3533_/CLK _3533_/D _3027_/Y vssd1 vssd1 vccd1 vccd1 _3533_/Q sky130_fd_sc_hd__dfrtp_1
Xhold815 _3477_/Q vssd1 vssd1 vccd1 vccd1 _2232_/A sky130_fd_sc_hd__buf_1
Xhold826 _2236_/X vssd1 vssd1 vccd1 vccd1 _3475_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold837 _1828_/X vssd1 vssd1 vccd1 vccd1 _3546_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold804 _3501_/Q vssd1 vssd1 vccd1 vccd1 hold804/X sky130_fd_sc_hd__dlygate4sd3_1
X_3464_ _3575_/CLK _3464_/D _2958_/Y vssd1 vssd1 vccd1 vccd1 _3464_/Q sky130_fd_sc_hd__dfrtp_1
Xhold859 _2253_/X vssd1 vssd1 vccd1 vccd1 _3468_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 _3150_/Q vssd1 vssd1 vccd1 vccd1 _1825_/A sky130_fd_sc_hd__clkbuf_2
X_2415_ _3580_/Q _2558_/B _2412_/X _2414_/Y vssd1 vssd1 vccd1 vccd1 _2415_/X sky130_fd_sc_hd__o211a_1
X_3395_ _3431_/CLK _3395_/D vssd1 vssd1 vccd1 vccd1 _3395_/Q sky130_fd_sc_hd__dfxtp_1
X_2346_ _1575_/Y _2208_/A _2205_/A _1576_/Y vssd1 vssd1 vccd1 vccd1 _2346_/X sky130_fd_sc_hd__o22a_1
X_2277_ _2271_/B _2281_/B _2271_/A vssd1 vssd1 vccd1 vccd1 _2278_/C sky130_fd_sc_hd__a21oi_1
Xclkbuf_2_2__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_2__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_15_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2023__B _2144_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2786__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xuart_macro_wrapper_133 vssd1 vssd1 vccd1 vccd1 uart_macro_wrapper_133/HI wbs_dat_o[22]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_80_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _2205_/A _2205_/B vssd1 vssd1 vccd1 vccd1 _2210_/C sky130_fd_sc_hd__nand2_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2710__A0 _2801_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3180_ _3413_/CLK _3180_/D vssd1 vssd1 vccd1 vccd1 _3180_/Q sky130_fd_sc_hd__dfxtp_1
X_2131_ _2146_/A _2381_/D vssd1 vssd1 vccd1 vccd1 _2133_/C sky130_fd_sc_hd__nand2_1
X_2062_ _3622_/Q _2070_/A vssd1 vssd1 vccd1 vccd1 _2064_/B sky130_fd_sc_hd__and2_2
XANTENNA__2823__S _2829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2964_ _3069_/A vssd1 vssd1 vccd1 vccd1 _2964_/Y sky130_fd_sc_hd__inv_2
X_1915_ _1912_/B _1918_/B _2546_/S vssd1 vssd1 vccd1 vccd1 _1916_/B sky130_fd_sc_hd__a21oi_1
X_2895_ hold642/X _2101_/Y _2900_/S vssd1 vssd1 vccd1 vccd1 _2895_/X sky130_fd_sc_hd__mux2_1
X_1846_ _1871_/A _1871_/B vssd1 vssd1 vccd1 vccd1 _1846_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold601 _2834_/X vssd1 vssd1 vccd1 vccd1 _3365_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold612 _3155_/Q vssd1 vssd1 vccd1 vccd1 hold612/X sky130_fd_sc_hd__dlygate4sd3_1
X_1777_ _3623_/Q _3622_/Q _1777_/C vssd1 vssd1 vccd1 vccd1 _2096_/A sky130_fd_sc_hd__or3_2
Xhold645 _2833_/X vssd1 vssd1 vccd1 vccd1 _3364_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 _3180_/Q vssd1 vssd1 vccd1 vccd1 hold634/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 _2626_/X vssd1 vssd1 vccd1 vccd1 _3173_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3516_ _3516_/CLK _3516_/D _3010_/Y vssd1 vssd1 vccd1 vccd1 _3516_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout101_A hold30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold656 _3408_/Q vssd1 vssd1 vccd1 vccd1 hold656/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 _2641_/X vssd1 vssd1 vccd1 vccd1 _3187_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold678 _3409_/Q vssd1 vssd1 vccd1 vccd1 hold678/X sky130_fd_sc_hd__dlygate4sd3_1
X_3447_ _3532_/CLK _3447_/D _2941_/Y vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__dfrtp_1
Xhold689 _2879_/X vssd1 vssd1 vccd1 vccd1 _3410_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ _3429_/CLK _3378_/D vssd1 vssd1 vccd1 vccd1 _3378_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2701__A0 _2803_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2329_ _3439_/Q _1598_/Y _2152_/B _2328_/X vssd1 vssd1 vccd1 vccd1 _2329_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_79_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2768__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1700_ _1700_/A _1700_/B vssd1 vssd1 vccd1 vccd1 _1700_/Y sky130_fd_sc_hd__nand2_1
X_2680_ _2802_/A1 hold163/X _2687_/S vssd1 vssd1 vccd1 vccd1 _2680_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1631_ hold80/X hold78/X hold12/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__mux2_1
XFILLER_0_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1562_ hold72/X vssd1 vssd1 vccd1 vccd1 _2325_/B sky130_fd_sc_hd__inv_2
X_3301_ _3319_/CLK _3301_/D vssd1 vssd1 vccd1 vccd1 _3301_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ _3509_/CLK _3232_/D vssd1 vssd1 vccd1 vccd1 _3232_/Q sky130_fd_sc_hd__dfxtp_1
X_3163_ _3438_/CLK _3163_/D vssd1 vssd1 vccd1 vccd1 _3163_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2114_ hold72/X _2383_/B vssd1 vssd1 vccd1 vccd1 _2116_/C sky130_fd_sc_hd__and2_1
X_3094_ _3124_/A vssd1 vssd1 vccd1 vccd1 _3094_/Y sky130_fd_sc_hd__inv_2
X_2045_ _3253_/Q _3130_/Q _3235_/Q _3226_/Q _2045_/S0 _2045_/S1 vssd1 vssd1 vccd1
+ vccd1 _2046_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1670__A0 _2400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2947_ _3122_/A vssd1 vssd1 vccd1 vccd1 _2947_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_72_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2878_ _2357_/B hold678/X _2880_/S vssd1 vssd1 vccd1 vccd1 _2878_/X sky130_fd_sc_hd__mux2_1
X_1829_ hold802/X _3545_/Q _1835_/S vssd1 vssd1 vccd1 vccd1 _1829_/X sky130_fd_sc_hd__mux2_1
Xhold420 _2245_/X vssd1 vssd1 vccd1 vccd1 _3472_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 _3482_/Q vssd1 vssd1 vccd1 vccd1 _2208_/A sky130_fd_sc_hd__clkbuf_2
Xhold442 _2662_/X vssd1 vssd1 vccd1 vccd1 _3203_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 _3221_/Q vssd1 vssd1 vccd1 vccd1 hold431/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 _2217_/X vssd1 vssd1 vccd1 vccd1 _3479_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 _2163_/X vssd1 vssd1 vccd1 vccd1 _3491_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 _3588_/Q vssd1 vssd1 vccd1 vccd1 _2334_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold497 _2824_/X vssd1 vssd1 vccd1 vccd1 _3356_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2728__S _2728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1632__S hold12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2801_ hold278/X _2801_/A1 _2809_/S vssd1 vssd1 vccd1 vccd1 _2801_/X sky130_fd_sc_hd__mux2_1
X_2732_ hold133/X _2802_/A1 _2739_/S vssd1 vssd1 vccd1 vccd1 _2732_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2663_ _2806_/A1 hold439/X _2666_/S vssd1 vssd1 vccd1 vccd1 _2663_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2904__A0 _2109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2594_ _2098_/S hold698/X _2601_/S vssd1 vssd1 vccd1 vccd1 _2594_/X sky130_fd_sc_hd__mux2_1
X_1614_ hold19/X hold51/X vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__nor2_1
XANTENNA__2402__A hold75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3215_ _3333_/CLK _3215_/D vssd1 vssd1 vccd1 vccd1 _3215_/Q sky130_fd_sc_hd__dfxtp_1
X_3146_ _3434_/CLK _3146_/D vssd1 vssd1 vccd1 vccd1 _3146_/Q sky130_fd_sc_hd__dfxtp_1
X_3077_ _3090_/A vssd1 vssd1 vccd1 vccd1 _3077_/Y sky130_fd_sc_hd__inv_2
X_2028_ _3246_/Q _3318_/Q _3309_/Q _3300_/Q _2049_/S0 _2219_/A vssd1 vssd1 vccd1 vccd1
+ _2028_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_9_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold250 _2715_/X vssd1 vssd1 vccd1 vccd1 _3249_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 _3217_/Q vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 input7/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 _2756_/X vssd1 vssd1 vccd1 vccd1 _3285_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 _2736_/X vssd1 vssd1 vccd1 vccd1 _3267_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2037__S1 _2219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 input7/A vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
X_3000_ _3101_/A vssd1 vssd1 vccd1 vccd1 _3000_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_52_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold87_A hold87/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2715_ _2806_/A1 hold249/X _2718_/S vssd1 vssd1 vccd1 vccd1 _2715_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2646_ _2358_/B hold770/X _2654_/S vssd1 vssd1 vccd1 vccd1 _2646_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2028__S1 _2219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2577_ hold1018/X _2577_/B vssd1 vssd1 vccd1 vccd1 _3577_/D sky130_fd_sc_hd__and2b_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3129_ _3129_/A vssd1 vssd1 vccd1 vccd1 _3129_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2741__S _2749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1919__A1 _1912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2003__A_N _2036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2977__A _3124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1759__C _1769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2651__S _2654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3480_ _3605_/CLK _3480_/D _2974_/Y vssd1 vssd1 vccd1 vccd1 _3480_/Q sky130_fd_sc_hd__dfrtp_1
X_2500_ _3186_/Q _3339_/Q _3168_/Q _3144_/Q _1944_/B _1943_/A vssd1 vssd1 vccd1 vccd1
+ _2500_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2583__A1 _2803_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2431_ _3172_/Q _3421_/Q _3412_/Q _3154_/Q _1918_/B _1912_/B vssd1 vssd1 vccd1 vccd1
+ _2431_/X sky130_fd_sc_hd__mux4_1
X_2362_ _1570_/Y _2098_/S _2109_/B _1569_/Y _2361_/X vssd1 vssd1 vccd1 vccd1 _2362_/X
+ sky130_fd_sc_hd__a221o_1
X_2293_ _3452_/Q hold15/X hold22/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__mux2_1
XANTENNA__2430__S1 _1912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2098__S _2098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_1__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2826__S _2829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2497__S1 _3518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_19_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3600_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2629_ _2103_/Y hold564/X _2633_/S vssd1 vssd1 vccd1 vccd1 _2629_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1640__S hold12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2646__S _2654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2980_ _3097_/A vssd1 vssd1 vccd1 vccd1 _2980_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_56_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1931_ _1931_/A _1931_/B vssd1 vssd1 vccd1 vccd1 _1934_/B sky130_fd_sc_hd__and2_1
X_1862_ _1861_/Y _1859_/B _1851_/A _1836_/A vssd1 vssd1 vccd1 vccd1 _1862_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_56_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput21 hold4/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__clkbuf_1
X_3601_ _3633_/CLK hold66/X _3092_/Y vssd1 vssd1 vccd1 vccd1 _3601_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput10 hold91/X vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput32 hold86/X vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__buf_1
X_1793_ _2387_/C _1793_/B vssd1 vssd1 vccd1 vccd1 _1793_/Y sky130_fd_sc_hd__nand2_1
Xhold816 _2231_/Y vssd1 vssd1 vccd1 vccd1 _3477_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3532_ _3532_/CLK _3532_/D _3026_/Y vssd1 vssd1 vccd1 vccd1 _3532_/Q sky130_fd_sc_hd__dfrtp_1
Xhold827 _3541_/Q vssd1 vssd1 vccd1 vccd1 hold827/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold805 _2055_/X vssd1 vssd1 vccd1 vccd1 _3501_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3463_ _3575_/CLK _3463_/D _2957_/Y vssd1 vssd1 vccd1 vccd1 _3463_/Q sky130_fd_sc_hd__dfrtp_1
Xhold838 _3544_/Q vssd1 vssd1 vccd1 vccd1 hold838/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 _1835_/S vssd1 vssd1 vccd1 vccd1 _1833_/S sky130_fd_sc_hd__clkbuf_2
X_2414_ _1578_/Y _2437_/A _2437_/B _2177_/A vssd1 vssd1 vccd1 vccd1 _2414_/Y sky130_fd_sc_hd__a22oi_1
X_3394_ _3438_/CLK _3394_/D vssd1 vssd1 vccd1 vccd1 _3394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2345_ _1576_/Y _2205_/A _2202_/A _1577_/Y _2344_/X vssd1 vssd1 vccd1 vccd1 _2345_/X
+ sky130_fd_sc_hd__a221o_1
X_2276_ _2272_/A _2278_/B _2275_/Y vssd1 vssd1 vccd1 vccd1 _2276_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2795__A1 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1635__S hold12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuart_macro_wrapper_134 vssd1 vssd1 vccd1 vccd1 uart_macro_wrapper_134/HI wbs_dat_o[24]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_21_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2130_ _2130_/A _2130_/B _2155_/B vssd1 vssd1 vccd1 vccd1 _2381_/D sky130_fd_sc_hd__or3_1
X_2061_ _2092_/A _2059_/Y _2060_/Y _2070_/A vssd1 vssd1 vccd1 vccd1 _2061_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2963_ _3069_/A vssd1 vssd1 vccd1 vccd1 _2963_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_56_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1914_ _1913_/A hold471/X _1911_/Y _2159_/B vssd1 vssd1 vccd1 vccd1 _3518_/D sky130_fd_sc_hd__a22o_1
XANTENNA__2405__A hold45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2777__A1 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2894_ hold518/X _2108_/Y _2900_/S vssd1 vssd1 vccd1 vccd1 _2894_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1845_ _1845_/A _1845_/B vssd1 vssd1 vccd1 vccd1 _1871_/B sky130_fd_sc_hd__and2_1
XFILLER_0_8_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold602 _3418_/Q vssd1 vssd1 vccd1 vccd1 hold602/X sky130_fd_sc_hd__dlygate4sd3_1
X_1776_ _3622_/Q _2070_/A vssd1 vssd1 vccd1 vccd1 _2065_/A sky130_fd_sc_hd__or2_1
XFILLER_0_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold635 _2633_/X vssd1 vssd1 vccd1 vccd1 _3180_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold613 _2605_/X vssd1 vssd1 vccd1 vccd1 _3155_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold624 _3145_/Q vssd1 vssd1 vccd1 vccd1 hold624/X sky130_fd_sc_hd__dlygate4sd3_1
X_3515_ _3516_/CLK _3515_/D _3009_/Y vssd1 vssd1 vccd1 vccd1 _3515_/Q sky130_fd_sc_hd__dfrtp_1
Xhold668 _3147_/Q vssd1 vssd1 vccd1 vccd1 hold668/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 _3407_/Q vssd1 vssd1 vccd1 vccd1 hold646/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 _2877_/X vssd1 vssd1 vccd1 vccd1 _3408_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 _2878_/X vssd1 vssd1 vccd1 vccd1 _3409_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3446_ _3589_/CLK _3446_/D _2940_/Y vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__dfrtp_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ _3429_/CLK _3377_/D vssd1 vssd1 vccd1 vccd1 _3377_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2328_ hold804/X _3349_/Q _1957_/B _3351_/Q _3348_/Q vssd1 vssd1 vccd1 vccd1 _2328_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2259_ _2259_/A _2259_/B _3473_/Q _2259_/D vssd1 vssd1 vccd1 vccd1 _2259_/X sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_34_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3571_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2759__A1 hold30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1630_ _3632_/Q hold15/X hold12/X vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__mux2_1
XFILLER_0_34_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3300_ _3318_/CLK _3300_/D vssd1 vssd1 vccd1 vccd1 _3300_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3056__A _3057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1561_ _3627_/Q vssd1 vssd1 vccd1 vccd1 _2116_/A sky130_fd_sc_hd__inv_2
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _3326_/CLK _3231_/D vssd1 vssd1 vccd1 vccd1 _3231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3162_ _3424_/CLK _3162_/D vssd1 vssd1 vccd1 vccd1 _3162_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2113_ _3627_/Q hold72/X _2113_/C hold99/X vssd1 vssd1 vccd1 vccd1 _2113_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_55_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3093_ _3101_/A vssd1 vssd1 vccd1 vccd1 _3093_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2044_ _2053_/A _2043_/Y _2055_/S vssd1 vssd1 vccd1 vccd1 _2044_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2542__S0 _1918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2946_ _3122_/A vssd1 vssd1 vccd1 vccd1 _2946_/Y sky130_fd_sc_hd__inv_2
X_2877_ _2360_/B hold656/X _2880_/S vssd1 vssd1 vccd1 vccd1 _2877_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1828_ hold836/X hold802/X _1835_/S vssd1 vssd1 vccd1 vccd1 _1828_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold410 _2589_/X vssd1 vssd1 vccd1 vccd1 _3138_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 _2212_/X vssd1 vssd1 vccd1 vccd1 _3482_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1759_ _1811_/S _3559_/Q _1769_/B vssd1 vssd1 vccd1 vccd1 _1759_/X sky130_fd_sc_hd__or3_1
Xhold421 _3241_/Q vssd1 vssd1 vccd1 vccd1 hold421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 _2683_/X vssd1 vssd1 vccd1 vccd1 _3221_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 _3329_/Q vssd1 vssd1 vccd1 vccd1 hold443/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 hold465/A vssd1 vssd1 vccd1 vccd1 _3579_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 _3518_/Q vssd1 vssd1 vccd1 vccd1 _1913_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold487 _2334_/Y vssd1 vssd1 vccd1 vccd1 _3382_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3429_ _3429_/CLK _3429_/D vssd1 vssd1 vccd1 vccd1 _3429_/Q sky130_fd_sc_hd__dfxtp_1
Xhold498 _3427_/Q vssd1 vssd1 vccd1 vccd1 hold498/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2686__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2744__S _2749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2610__A0 _2357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2654__S _2654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1652__A1 _2400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2800_ _2800_/A _2800_/B vssd1 vssd1 vccd1 vccd1 _2809_/S sky130_fd_sc_hd__nor2_4
X_2731_ hold224/X _2801_/A1 _2739_/S vssd1 vssd1 vccd1 vccd1 _2731_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2601__A0 _2356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2662_ _2805_/A1 hold441/X _2666_/S vssd1 vssd1 vccd1 vccd1 _2662_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2593_ _2358_/B hold594/X _2601_/S vssd1 vssd1 vccd1 vccd1 _2593_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1613_ hold92/A hold50/X _1623_/C hold8/X vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__or4bb_1
XANTENNA__2829__S _2829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3214_ _3509_/CLK _3214_/D vssd1 vssd1 vccd1 vccd1 _3214_/Q sky130_fd_sc_hd__dfxtp_1
X_3145_ _3521_/CLK _3145_/D vssd1 vssd1 vccd1 vccd1 _3145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3076_ _3090_/A vssd1 vssd1 vccd1 vccd1 _3076_/Y sky130_fd_sc_hd__inv_2
X_2027_ _3291_/Q _3282_/Q _3273_/Q _3264_/Q _2221_/B _2219_/A vssd1 vssd1 vccd1 vccd1
+ _2027_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2515__S0 _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2929_ _3127_/A vssd1 vssd1 vccd1 vccd1 _2929_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_60_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold240 _2778_/X vssd1 vssd1 vccd1 vccd1 _3305_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 _3323_/Q vssd1 vssd1 vccd1 vccd1 hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _2679_/X vssd1 vssd1 vccd1 vccd1 _3217_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _3276_/Q vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 _1674_/C vssd1 vssd1 vccd1 vccd1 _1659_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 _3248_/Q vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2659__A0 _2802_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout74_A _2103_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1634__A1 _2406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2831__A0 _2358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2649__S _2654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2362__A2 _2098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 input8/A vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_0__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_3_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2714_ _2805_/A1 hold284/X _2718_/S vssd1 vssd1 vccd1 vccd1 _2714_/X sky130_fd_sc_hd__mux2_1
X_2645_ _2901_/A _2830_/B vssd1 vssd1 vccd1 vccd1 _2654_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_42_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2576_ _2576_/A hold98/X _2576_/C vssd1 vssd1 vccd1 vccd1 _2576_/X sky130_fd_sc_hd__and3_1
X_3128_ _3129_/A vssd1 vssd1 vccd1 vccd1 _3128_/Y sky130_fd_sc_hd__inv_2
X_3059_ _3061_/A vssd1 vssd1 vccd1 vccd1 _3059_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1919__A2 _1918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1638__S hold12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2042__B _2144_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2469__S _3518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2032__A1 _2144_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2430_ _3371_/Q _3353_/Q _3362_/Q _3190_/Q _1918_/B _1912_/B vssd1 vssd1 vccd1 vccd1
+ _2430_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2335__A2 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2361_ _1567_/Y _2104_/B _2359_/X _2360_/Y vssd1 vssd1 vccd1 vccd1 _2361_/X sky130_fd_sc_hd__a2bb2o_1
X_2292_ _3453_/Q hold25/X hold22/X vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__mux2_1
XFILLER_0_47_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2842__S _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout124_A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_2_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2628_ _2105_/A hold706/X _2633_/S vssd1 vssd1 vccd1 vccd1 _2628_/X sky130_fd_sc_hd__mux2_1
X_2559_ _2572_/C _2559_/B _2572_/D vssd1 vssd1 vccd1 vccd1 _2559_/X sky130_fd_sc_hd__and3_1
XFILLER_0_84_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1930_ _1934_/A _1930_/B vssd1 vssd1 vccd1 vccd1 _1931_/B sky130_fd_sc_hd__nor2_1
X_1861_ _1851_/A _1851_/B _1837_/A vssd1 vssd1 vccd1 vccd1 _1861_/Y sky130_fd_sc_hd__o21ai_1
Xinput22 hold77/X vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__clkbuf_2
Xinput11 hold7/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__buf_1
X_3600_ _3600_/CLK _3600_/D _3091_/Y vssd1 vssd1 vccd1 vccd1 _3600_/Q sky130_fd_sc_hd__dfrtp_1
X_3531_ _3532_/CLK _3531_/D _3025_/Y vssd1 vssd1 vccd1 vccd1 _3531_/Q sky130_fd_sc_hd__dfrtp_1
X_1792_ _1792_/A _1792_/B _1792_/C _1792_/D vssd1 vssd1 vccd1 vccd1 _1793_/B sky130_fd_sc_hd__and4_1
Xinput33 hold44/X vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__clkbuf_1
Xhold806 _3461_/Q vssd1 vssd1 vccd1 vccd1 hold806/X sky130_fd_sc_hd__buf_1
Xhold817 _3515_/Q vssd1 vssd1 vccd1 vccd1 hold817/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 _1834_/X vssd1 vssd1 vccd1 vccd1 _3540_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3462_ _3574_/CLK _3462_/D _2956_/Y vssd1 vssd1 vccd1 vccd1 _3462_/Q sky130_fd_sc_hd__dfrtp_4
Xhold839 _1831_/X vssd1 vssd1 vccd1 vccd1 _3543_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3393_ _3438_/CLK _3393_/D vssd1 vssd1 vccd1 vccd1 _3393_/Q sky130_fd_sc_hd__dfxtp_1
X_2413_ _2413_/A _2413_/B vssd1 vssd1 vccd1 vccd1 _2437_/B sky130_fd_sc_hd__nor2_1
X_2344_ _1577_/Y _2202_/A _2217_/S _1578_/Y vssd1 vssd1 vccd1 vccd1 _2344_/X sky130_fd_sc_hd__o22a_1
X_2275_ _2283_/A _2275_/B vssd1 vssd1 vccd1 vccd1 _2275_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2747__S _2749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2482__S _2546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xuart_macro_wrapper_135 vssd1 vssd1 vccd1 vccd1 uart_macro_wrapper_135/HI wbs_dat_o[29]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_4_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3610_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2060_ _3547_/Q _2084_/B _2092_/A vssd1 vssd1 vccd1 vccd1 _2060_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2962_ _3069_/A vssd1 vssd1 vccd1 vccd1 _2962_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1913_ _1913_/A _1916_/A vssd1 vssd1 vccd1 vccd1 _2159_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_29_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2893_ hold530/X _2087_/Y _2900_/S vssd1 vssd1 vccd1 vccd1 _2893_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1844_ _1845_/B vssd1 vssd1 vccd1 vccd1 _1844_/Y sky130_fd_sc_hd__inv_2
Xhold603 _2888_/X vssd1 vssd1 vccd1 vccd1 _3418_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1775_ _3622_/Q _2070_/A vssd1 vssd1 vccd1 vccd1 _2064_/A sky130_fd_sc_hd__nor2_4
XANTENNA_hold62_A hold62/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold614 _3395_/Q vssd1 vssd1 vccd1 vccd1 hold614/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 _2599_/X vssd1 vssd1 vccd1 vccd1 _3145_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 _3367_/Q vssd1 vssd1 vccd1 vccd1 hold636/X sky130_fd_sc_hd__dlygate4sd3_1
X_3514_ _3602_/CLK _3514_/D _3008_/Y vssd1 vssd1 vccd1 vccd1 _3514_/Q sky130_fd_sc_hd__dfrtp_1
X_3445_ _3589_/CLK _3445_/D _2939_/Y vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__dfrtp_1
Xhold658 _3378_/Q vssd1 vssd1 vccd1 vccd1 hold658/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 _2876_/X vssd1 vssd1 vccd1 vccd1 _3407_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold669 _2601_/X vssd1 vssd1 vccd1 vccd1 _3147_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _3516_/CLK _3376_/D vssd1 vssd1 vccd1 vccd1 _3376_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2327_ _2326_/X hold99/X _2116_/A _2325_/X vssd1 vssd1 vccd1 vccd1 _2327_/X sky130_fd_sc_hd__a2bb2o_1
X_2258_ _3463_/Q hold778/X _3462_/Q vssd1 vssd1 vccd1 vccd1 _2258_/X sky130_fd_sc_hd__mux2_1
X_2189_ _2186_/X _2241_/B _2225_/A _2193_/B vssd1 vssd1 vccd1 vccd1 _3486_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1560_ _1560_/A vssd1 vssd1 vccd1 vccd1 _2550_/A sky130_fd_sc_hd__inv_2
XFILLER_0_22_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _3326_/CLK _3230_/D vssd1 vssd1 vccd1 vccd1 _3230_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ _3579_/CLK _3161_/D vssd1 vssd1 vccd1 vccd1 _3161_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2695__A1 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2112_ _3627_/Q hold99/X _2325_/B _2113_/C vssd1 vssd1 vccd1 vccd1 _2112_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_55_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3092_ _3122_/A vssd1 vssd1 vccd1 vccd1 _3092_/Y sky130_fd_sc_hd__inv_2
X_2043_ _2144_/C _2041_/Y _2042_/Y vssd1 vssd1 vccd1 vccd1 _2043_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2542__S1 _1912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2945_ _3122_/A vssd1 vssd1 vccd1 vccd1 _2945_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2135__B _2144_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2876_ _2104_/B hold646/X _2880_/S vssd1 vssd1 vccd1 vccd1 _2876_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1827_ _2383_/B hold836/X _1833_/S vssd1 vssd1 vccd1 vccd1 _3547_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold411 _3223_/Q vssd1 vssd1 vccd1 vccd1 hold411/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold400 _2666_/X vssd1 vssd1 vccd1 vccd1 _3207_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1758_ _1755_/B _2387_/C _1757_/X vssd1 vssd1 vccd1 vccd1 _1758_/X sky130_fd_sc_hd__o21a_1
Xhold422 _2705_/X vssd1 vssd1 vccd1 vccd1 _3241_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 _3216_/Q vssd1 vssd1 vccd1 vccd1 hold433/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 _2805_/X vssd1 vssd1 vccd1 vccd1 _3329_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold455 _3480_/Q vssd1 vssd1 vccd1 vccd1 _2202_/A sky130_fd_sc_hd__clkbuf_2
X_1689_ _1689_/A _1689_/B _1708_/B vssd1 vssd1 vccd1 vccd1 _1704_/B sky130_fd_sc_hd__or3_1
Xhold477 _3517_/Q vssd1 vssd1 vccd1 vccd1 hold477/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 hold466/A vssd1 vssd1 vccd1 vccd1 _1935_/A sky130_fd_sc_hd__buf_2
X_3428_ _3579_/CLK _3428_/D vssd1 vssd1 vccd1 vccd1 _3428_/Q sky130_fd_sc_hd__dfxtp_1
Xhold488 _3360_/Q vssd1 vssd1 vccd1 vccd1 hold488/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold499 _2898_/X vssd1 vssd1 vccd1 vccd1 _3427_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3359_ _3429_/CLK _3359_/D vssd1 vssd1 vccd1 vccd1 _3359_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2000__S _2000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2361__A2_N _2104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2730_ _2800_/A _2760_/B vssd1 vssd1 vccd1 vccd1 _2739_/S sky130_fd_sc_hd__nor2_4
X_2661_ _2804_/A1 hold210/X _2666_/S vssd1 vssd1 vccd1 vccd1 _2661_/X sky130_fd_sc_hd__mux2_1
X_1612_ _1612_/A _1612_/B _1624_/B hold18/X vssd1 vssd1 vccd1 vccd1 _1612_/X sky130_fd_sc_hd__or4_1
X_2592_ _2810_/B _2901_/A vssd1 vssd1 vccd1 vccd1 _2601_/S sky130_fd_sc_hd__nand2_4
XANTENNA__2365__B1 _2103_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2117__B1 _1769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3213_ _3330_/CLK _3213_/D vssd1 vssd1 vccd1 vccd1 _3213_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2668__A1 _2801_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3144_ _3408_/CLK _3144_/D vssd1 vssd1 vccd1 vccd1 _3144_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2845__S _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3075_ _3090_/A vssd1 vssd1 vccd1 vccd1 _3075_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2515__S1 _1943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2026_ _3219_/Q _3210_/Q _3201_/Q _3327_/Q _2045_/S0 _2195_/A1 vssd1 vssd1 vccd1
+ vccd1 _2026_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_49_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2928_ _3127_/A vssd1 vssd1 vccd1 vccd1 _2928_/Y sky130_fd_sc_hd__inv_2
X_2859_ _2355_/B hold652/X _2860_/S vssd1 vssd1 vccd1 vccd1 _2859_/X sky130_fd_sc_hd__mux2_1
Xhold252 _2798_/X vssd1 vssd1 vccd1 vccd1 _3323_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 _3211_/Q vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 _3332_/Q vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 _3312_/Q vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _2746_/X vssd1 vssd1 vccd1 vccd1 _3276_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 _2575_/X vssd1 vssd1 vccd1 vccd1 _3602_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 _2714_/X vssd1 vssd1 vccd1 vccd1 _3248_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2595__A0 _2109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput9 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_59_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2822__A1 _2098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2713_ _2804_/A1 hold157/X _2718_/S vssd1 vssd1 vccd1 vccd1 _2713_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2644_ _3522_/Q _3521_/Q vssd1 vssd1 vccd1 vccd1 _2830_/B sky130_fd_sc_hd__and2b_2
X_2575_ _2576_/A hold98/A _2575_/C vssd1 vssd1 vccd1 vccd1 _2575_/X sky130_fd_sc_hd__and3_1
XFILLER_0_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3127_ _3127_/A vssd1 vssd1 vccd1 vccd1 _3127_/Y sky130_fd_sc_hd__inv_2
X_3058_ _3061_/A vssd1 vssd1 vccd1 vccd1 _3058_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2813__A1 _2109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2009_ _2315_/A1 _2007_/X _2008_/Y _2003_/Y vssd1 vssd1 vccd1 vccd1 _2009_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2485__S _3517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2804__A1 _2804_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2360_ _3616_/Q _2360_/B vssd1 vssd1 vccd1 vccd1 _2360_/Y sky130_fd_sc_hd__nand2_1
X_2291_ _3454_/Q hold2/X hold22/A vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__mux2_1
XFILLER_0_2_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold92_A hold92/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout117_A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2627_ _2109_/B hold752/X _2633_/S vssd1 vssd1 vccd1 vccd1 _2627_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_28_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3550_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2558_ hold64/A _2558_/B _2558_/C vssd1 vssd1 vccd1 vccd1 _2572_/D sky130_fd_sc_hd__and3_1
XFILLER_0_2_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2489_ _3584_/Q hold95/A _2410_/X _3346_/Q _2488_/X vssd1 vssd1 vccd1 vccd1 _2489_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2053__B _2144_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2722__A0 _2803_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2789__A0 hold30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1860_ _1837_/A _1852_/Y _1859_/X _1859_/A _1836_/A vssd1 vssd1 vccd1 vccd1 _1860_/X
+ sky130_fd_sc_hd__a32o_1
Xinput12 input12/A vssd1 vssd1 vccd1 vccd1 _1623_/C sky130_fd_sc_hd__clkbuf_2
X_1791_ _1791_/A _2126_/B vssd1 vssd1 vccd1 vccd1 _1792_/D sky130_fd_sc_hd__nand2_1
X_3530_ _3532_/CLK _3530_/D _3024_/Y vssd1 vssd1 vccd1 vccd1 _3530_/Q sky130_fd_sc_hd__dfrtp_1
Xinput34 hold29/X vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__buf_1
Xinput23 hold14/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__buf_1
Xhold807 _2274_/Y vssd1 vssd1 vccd1 vccd1 _3461_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold818 _3575_/Q vssd1 vssd1 vccd1 vccd1 _1697_/A sky130_fd_sc_hd__dlygate4sd3_1
X_3461_ _3594_/CLK _3461_/D _2955_/Y vssd1 vssd1 vccd1 vccd1 _3461_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold829 _3574_/Q vssd1 vssd1 vccd1 vccd1 _1697_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2713__A0 _2804_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3392_ _3521_/CLK _3392_/D vssd1 vssd1 vccd1 vccd1 _3392_/Q sky130_fd_sc_hd__dfxtp_1
X_2412_ _3592_/Q _2438_/B _2558_/C _3590_/Q vssd1 vssd1 vccd1 vccd1 _2412_/X sky130_fd_sc_hd__o22a_1
X_2343_ _2343_/A _2343_/B vssd1 vssd1 vccd1 vccd1 _2343_/Y sky130_fd_sc_hd__nor2_1
X_2274_ hold806/X _2275_/B _2273_/Y vssd1 vssd1 vccd1 vccd1 _2274_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1989_ hold788/X _1988_/Y _2000_/S vssd1 vssd1 vccd1 vccd1 _1989_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2704__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2763__S _2769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2064__A _2064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuart_macro_wrapper_136 vssd1 vssd1 vccd1 vccd1 io_oeb[0] uart_macro_wrapper_136/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_2_3__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2961_ _3069_/A vssd1 vssd1 vccd1 vccd1 _2961_/Y sky130_fd_sc_hd__inv_2
X_1912_ _2546_/S _1912_/B _1918_/B vssd1 vssd1 vccd1 vccd1 _1916_/A sky130_fd_sc_hd__and3_1
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2892_ hold538/X _2097_/X _2900_/S vssd1 vssd1 vccd1 vccd1 _2892_/X sky130_fd_sc_hd__mux2_1
X_1843_ _1843_/A _1877_/A _1877_/B vssd1 vssd1 vccd1 vccd1 _1845_/B sky130_fd_sc_hd__and3_1
X_1774_ _3623_/Q _3622_/Q vssd1 vssd1 vccd1 vccd1 _1774_/X sky130_fd_sc_hd__or2_1
Xhold626 _3172_/Q vssd1 vssd1 vccd1 vccd1 hold626/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold615 _2863_/X vssd1 vssd1 vccd1 vccd1 _3395_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold604 _3334_/Q vssd1 vssd1 vccd1 vccd1 hold604/X sky130_fd_sc_hd__dlygate4sd3_1
X_3513_ _3602_/CLK _3513_/D _3007_/Y vssd1 vssd1 vccd1 vccd1 _3513_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold659 _2848_/X vssd1 vssd1 vccd1 vccd1 _3378_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 _3179_/Q vssd1 vssd1 vccd1 vccd1 hold648/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold637 _2836_/X vssd1 vssd1 vccd1 vccd1 _3367_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3444_ _3635_/CLK _3444_/D _2938_/Y vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__2848__S _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ _3431_/CLK _3375_/D vssd1 vssd1 vccd1 vccd1 _3375_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2326_ _2116_/A _2325_/C _2325_/B vssd1 vssd1 vccd1 vccd1 _2326_/X sky130_fd_sc_hd__a21o_1
X_2257_ hold878/X hold898/X _3462_/Q vssd1 vssd1 vccd1 vccd1 _2257_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2583__S _2589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2188_ _2225_/A _2191_/A vssd1 vssd1 vccd1 vccd1 _2241_/B sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_43_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3619_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout97_A _3483_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _3575_/CLK _3160_/D vssd1 vssd1 vccd1 vccd1 _3160_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1 wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
X_2111_ _2111_/A _2111_/B vssd1 vssd1 vccd1 vccd1 _2113_/C sky130_fd_sc_hd__xnor2_1
X_3091_ input2/X vssd1 vssd1 vccd1 vccd1 _3091_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2042_ _3503_/Q _2144_/C vssd1 vssd1 vccd1 vccd1 _2042_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_69_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2944_ _3122_/A vssd1 vssd1 vccd1 vccd1 _2944_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1958__A1 _2144_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2875_ _2105_/A hold664/X _2880_/S vssd1 vssd1 vccd1 vccd1 _2875_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1826_ _1833_/S vssd1 vssd1 vccd1 vccd1 _1826_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2907__A0 _2360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold401 _3259_/Q vssd1 vssd1 vccd1 vccd1 hold401/X sky130_fd_sc_hd__dlygate4sd3_1
X_1757_ _1811_/S _1757_/B _1769_/B vssd1 vssd1 vccd1 vccd1 _1757_/X sky130_fd_sc_hd__or3_1
XFILLER_0_20_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold445 _3234_/Q vssd1 vssd1 vccd1 vccd1 hold445/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 _2685_/X vssd1 vssd1 vccd1 vccd1 _3223_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 _2676_/X vssd1 vssd1 vccd1 vccd1 _3216_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 _3130_/Q vssd1 vssd1 vccd1 vccd1 hold423/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold456 _2216_/X vssd1 vssd1 vccd1 vccd1 _3480_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 _3582_/Q vssd1 vssd1 vccd1 vccd1 hold478/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 _1919_/Y vssd1 vssd1 vccd1 vccd1 hold467/X sky130_fd_sc_hd__dlygate4sd3_1
X_1688_ _3590_/Q _3472_/Q hold840/X vssd1 vssd1 vccd1 vccd1 _1688_/X sky130_fd_sc_hd__o21ba_1
Xhold489 _2828_/X vssd1 vssd1 vccd1 vccd1 _3360_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3427_ _3575_/CLK _3427_/D vssd1 vssd1 vccd1 vccd1 _3427_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3358_ _3516_/CLK _3358_/D vssd1 vssd1 vccd1 vccd1 _3358_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2309_ _2309_/A _2309_/B vssd1 vssd1 vccd1 vccd1 _2310_/B sky130_fd_sc_hd__xnor2_1
X_3289_ _3324_/CLK _3289_/D vssd1 vssd1 vccd1 vccd1 _3289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2049__S1 _2195_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold990 _2234_/X vssd1 vssd1 vccd1 vccd1 _3476_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1980__S0 _2045_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2660_ _2803_/A1 hold355/X _2666_/S vssd1 vssd1 vccd1 vccd1 _2660_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1611_ hold34/X _1611_/B vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__nor2_2
XFILLER_0_41_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2591_ _3520_/Q _3519_/Q _2613_/B vssd1 vssd1 vccd1 vccd1 _2901_/A sky130_fd_sc_hd__and3_4
XFILLER_0_5_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3212_ _3329_/CLK _3212_/D vssd1 vssd1 vccd1 vccd1 _3212_/Q sky130_fd_sc_hd__dfxtp_1
X_3143_ _3433_/CLK _3143_/D vssd1 vssd1 vccd1 vccd1 _3143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3074_ _3101_/A vssd1 vssd1 vccd1 vccd1 _3074_/Y sky130_fd_sc_hd__inv_2
X_2025_ _2036_/S _2025_/B vssd1 vssd1 vccd1 vccd1 _2025_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2927_ _3129_/A vssd1 vssd1 vccd1 vccd1 _2927_/Y sky130_fd_sc_hd__inv_2
X_2858_ _2357_/B hold720/X _2860_/S vssd1 vssd1 vccd1 vccd1 _2858_/X sky130_fd_sc_hd__mux2_1
X_2789_ hold30/X _2789_/A1 hold38/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__mux2_1
Xhold220 _3244_/Q vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
X_1809_ _1809_/A _1809_/B vssd1 vssd1 vccd1 vccd1 _1810_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_13_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold242 _2671_/X vssd1 vssd1 vccd1 vccd1 _3211_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 _2808_/X vssd1 vssd1 vccd1 vccd1 _3332_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 _3226_/Q vssd1 vssd1 vccd1 vccd1 hold253/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 _3303_/Q vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _2786_/X vssd1 vssd1 vccd1 vccd1 _3312_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 _3592_/Q vssd1 vssd1 vccd1 vccd1 hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 _3275_/Q vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2771__S _2779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2712_ _2803_/A1 hold345/X _2718_/S vssd1 vssd1 vccd1 vccd1 _2712_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2586__A1 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2643_ _2356_/B hold578/X _2643_/S vssd1 vssd1 vccd1 vccd1 _2643_/X sky130_fd_sc_hd__mux2_1
X_2574_ _2574_/A hold21/A _2574_/C vssd1 vssd1 vccd1 vccd1 _3655_/A sky130_fd_sc_hd__and3_4
X_3126_ _3127_/A vssd1 vssd1 vccd1 vccd1 _3126_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3057_ _3057_/A vssd1 vssd1 vccd1 vccd1 _3057_/Y sky130_fd_sc_hd__inv_2
X_2008_ _2036_/S _2004_/X _2315_/A1 vssd1 vssd1 vccd1 vccd1 _2008_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_37_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2329__A1 _3439_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold476_A _3518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2766__S _2769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2290_ _3455_/Q hold56/X hold22/X vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__mux2_1
XANTENNA_output60_A _3655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2626_ _2098_/S hold622/X _2633_/S vssd1 vssd1 vccd1 vccd1 _2626_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2731__A1 _2801_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2557_ _3630_/Q hold11/A vssd1 vssd1 vccd1 vccd1 _2557_/X sky130_fd_sc_hd__or2_1
X_2488_ _3346_/Q _1675_/X _2409_/Y hold85/A vssd1 vssd1 vccd1 vccd1 _2488_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2586__S _2589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3109_ _3129_/A vssd1 vssd1 vccd1 vccd1 _3109_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2798__A1 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput13 input13/A vssd1 vssd1 vccd1 vccd1 _1612_/B sky130_fd_sc_hd__buf_1
X_1790_ _1791_/A _2126_/B vssd1 vssd1 vccd1 vccd1 _1792_/C sky130_fd_sc_hd__or2_1
Xinput24 hold24/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__clkbuf_1
Xinput35 hold58/X vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__buf_1
XFILLER_0_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold808 _3520_/Q vssd1 vssd1 vccd1 vccd1 _1902_/A sky130_fd_sc_hd__buf_1
Xhold819 _1694_/X vssd1 vssd1 vccd1 vccd1 _3575_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3460_ _3594_/CLK _3460_/D _2954_/Y vssd1 vssd1 vccd1 vccd1 _3460_/Q sky130_fd_sc_hd__dfrtp_1
X_3391_ _3521_/CLK _3391_/D vssd1 vssd1 vccd1 vccd1 _3391_/Q sky130_fd_sc_hd__dfxtp_1
X_2411_ _2165_/B hold20/A hold63/A vssd1 vssd1 vccd1 vccd1 _2558_/C sky130_fd_sc_hd__o21ai_4
X_2342_ _2339_/X _2340_/X _2341_/X _1595_/Y vssd1 vssd1 vccd1 vccd1 _2343_/B sky130_fd_sc_hd__o31a_1
X_2273_ hold806/X _2275_/B _2283_/A vssd1 vssd1 vccd1 vccd1 _2273_/Y sky130_fd_sc_hd__o21bai_1
XANTENNA__3091__A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1988_ _1988_/A vssd1 vssd1 vccd1 vccd1 _1988_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_70_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3589_ _3589_/CLK hold96/X _3080_/Y vssd1 vssd1 vccd1 vccd1 _3589_/Q sky130_fd_sc_hd__dfrtp_1
X_2609_ _2360_/B hold532/X _2612_/S vssd1 vssd1 vccd1 vccd1 _2609_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2640__A0 _2360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_88_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1682__A1 hold70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2960_ _3069_/A vssd1 vssd1 vccd1 vccd1 _2960_/Y sky130_fd_sc_hd__inv_2
X_2891_ _2891_/A _2891_/B vssd1 vssd1 vccd1 vccd1 _2900_/S sky130_fd_sc_hd__and2_4
XANTENNA__2631__A0 _2357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1911_ _1935_/A _1911_/B vssd1 vssd1 vccd1 vccd1 _1911_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1842_ _1877_/A _1877_/B vssd1 vssd1 vccd1 vccd1 _1842_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1773_ _2383_/A _1795_/B vssd1 vssd1 vccd1 vccd1 _1773_/Y sky130_fd_sc_hd__nor2_1
Xhold616 _3438_/Q vssd1 vssd1 vccd1 vccd1 hold616/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 _2625_/X vssd1 vssd1 vccd1 vccd1 _3172_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold605 _2811_/X vssd1 vssd1 vccd1 vccd1 _3334_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3512_ _3614_/CLK _3512_/D _3006_/Y vssd1 vssd1 vccd1 vccd1 _3512_/Q sky130_fd_sc_hd__dfrtp_1
Xhold649 _2632_/X vssd1 vssd1 vccd1 vccd1 _3179_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 _3417_/Q vssd1 vssd1 vccd1 vccd1 hold638/X sky130_fd_sc_hd__dlygate4sd3_1
X_3443_ _3635_/CLK _3443_/D _2937_/Y vssd1 vssd1 vccd1 vccd1 _3443_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _3413_/CLK _3374_/D vssd1 vssd1 vccd1 vccd1 _3374_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2325_ hold99/X _2325_/B _2325_/C vssd1 vssd1 vccd1 vccd1 _2325_/X sky130_fd_sc_hd__and3_1
X_2256_ _2249_/A hold878/X _3462_/Q vssd1 vssd1 vccd1 vccd1 _2256_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2864__S _2870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2545__S0 _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2187_ _2222_/A _2219_/A _2221_/B vssd1 vssd1 vccd1 vccd1 _2191_/A sky130_fd_sc_hd__and3_1
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2622__A0 _2355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3318_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2774__S _2779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1664__A1 _2399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2075__A _2356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
X_2110_ _2110_/A _2110_/B vssd1 vssd1 vccd1 vccd1 _2111_/B sky130_fd_sc_hd__xnor2_1
X_3090_ _3090_/A vssd1 vssd1 vccd1 vccd1 _3090_/Y sky130_fd_sc_hd__inv_2
X_2041_ _2315_/A1 _2036_/X _2040_/X vssd1 vssd1 vccd1 vccd1 _2041_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__2852__A0 _2358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2943_ _3032_/A vssd1 vssd1 vccd1 vccd1 _2943_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2604__A0 _2358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2874_ _2109_/B hold684/X _2880_/S vssd1 vssd1 vccd1 vccd1 _2874_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1825_ _1825_/A _2387_/C vssd1 vssd1 vccd1 vccd1 _1835_/S sky130_fd_sc_hd__nand2_4
X_1756_ _1753_/B _2387_/C _1755_/X vssd1 vssd1 vccd1 vccd1 _1756_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_4_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold402 _2726_/X vssd1 vssd1 vccd1 vccd1 _3259_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 _3136_/Q vssd1 vssd1 vccd1 vccd1 hold435/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 _3333_/Q vssd1 vssd1 vccd1 vccd1 hold413/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 _2581_/X vssd1 vssd1 vccd1 vccd1 _3130_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold457 _3481_/Q vssd1 vssd1 vccd1 vccd1 _2205_/A sky130_fd_sc_hd__clkbuf_2
X_1687_ hold275/X _2576_/A hold65/X vssd1 vssd1 vccd1 vccd1 _3592_/D sky130_fd_sc_hd__mux2_1
Xhold468 _1920_/X vssd1 vssd1 vccd1 vccd1 _3516_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 _2697_/X vssd1 vssd1 vccd1 vccd1 _3234_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold479 _2348_/Y vssd1 vssd1 vccd1 vccd1 _3345_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3426_ _3516_/CLK _3426_/D vssd1 vssd1 vccd1 vccd1 _3426_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3357_ _3431_/CLK _3357_/D vssd1 vssd1 vccd1 vccd1 _3357_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _1967_/B _2308_/B vssd1 vssd1 vccd1 vccd1 _2309_/B sky130_fd_sc_hd__and2b_1
X_3288_ _3484_/CLK hold43/X vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__2518__S0 _2532_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2239_ _2381_/B _2381_/C _2363_/A _1591_/Y vssd1 vssd1 vccd1 vccd1 _2239_/X sky130_fd_sc_hd__o31a_1
XANTENNA__1646__A1 _2406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2769__S _2769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold980 _1754_/X vssd1 vssd1 vccd1 vccd1 _3563_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold991 _3553_/Q vssd1 vssd1 vccd1 vccd1 _1771_/B sky130_fd_sc_hd__buf_1
XANTENNA__1980__S1 _2045_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2834__A0 _2101_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1637__A1 hold70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1610_ _1657_/A hold62/A input4/X input5/X vssd1 vssd1 vccd1 vccd1 _1610_/X sky130_fd_sc_hd__or4_1
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2590_ _3521_/Q _3522_/Q vssd1 vssd1 vccd1 vccd1 _2810_/B sky130_fd_sc_hd__and2b_2
XFILLER_0_22_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2365__A2 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3211_ _3509_/CLK _3211_/D vssd1 vssd1 vccd1 vccd1 _3211_/Q sky130_fd_sc_hd__dfxtp_1
X_3142_ _3433_/CLK _3142_/D vssd1 vssd1 vccd1 vccd1 _3142_/Q sky130_fd_sc_hd__dfxtp_1
X_3073_ _3097_/A vssd1 vssd1 vccd1 vccd1 _3073_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_82_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2024_ _3255_/Q _3132_/Q _3237_/Q _3228_/Q _2045_/S0 _2045_/S1 vssd1 vssd1 vccd1
+ vccd1 _2025_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_72_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2926_ _3054_/A vssd1 vssd1 vccd1 vccd1 _2926_/Y sky130_fd_sc_hd__inv_2
X_2857_ _2360_/B hold742/X _2860_/S vssd1 vssd1 vccd1 vccd1 _2857_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1808_ _1808_/A _1808_/B _1825_/A _1808_/D vssd1 vssd1 vccd1 vccd1 _1809_/B sky130_fd_sc_hd__or4_1
X_2788_ _2808_/A1 hold233/X hold38/X vssd1 vssd1 vccd1 vccd1 _2788_/X sky130_fd_sc_hd__mux2_1
Xhold210 _3202_/Q vssd1 vssd1 vccd1 vccd1 hold210/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 _2710_/X vssd1 vssd1 vccd1 vccd1 _3244_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1739_ _1739_/A _1739_/B _1739_/C _1739_/D vssd1 vssd1 vccd1 vccd1 _2381_/C sky130_fd_sc_hd__or4_2
XANTENNA__2589__S _2589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold232 _3621_/Q vssd1 vssd1 vccd1 vccd1 _1777_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 _3328_/Q vssd1 vssd1 vccd1 vccd1 hold243/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 _3316_/Q vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 _2776_/X vssd1 vssd1 vccd1 vccd1 _3303_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 _2689_/X vssd1 vssd1 vccd1 vccd1 _3226_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 _3266_/Q vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__dlygate4sd3_1
X_3409_ _3521_/CLK _3409_/D vssd1 vssd1 vccd1 vccd1 _3409_/Q sky130_fd_sc_hd__dfxtp_1
Xhold298 _2745_/X vssd1 vssd1 vccd1 vccd1 _3275_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1962__S1 _2195_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1619__A1 _2401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold888_A _2198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2711_ _2802_/A1 hold131/X _2718_/S vssd1 vssd1 vccd1 vccd1 _2711_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2642_ _2355_/B hold680/X _2643_/S vssd1 vssd1 vccd1 vccd1 _2642_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2573_ _3455_/Q hold21/A _2574_/C _2574_/A vssd1 vssd1 vccd1 vccd1 _2573_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3094__A _3124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1607__A _1607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold30_A hold30/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3125_ _3127_/A vssd1 vssd1 vccd1 vccd1 _3125_/Y sky130_fd_sc_hd__inv_2
X_3056_ _3057_/A vssd1 vssd1 vccd1 vccd1 _3056_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2872__S _2880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2007_ _2006_/X _2005_/X _2036_/S vssd1 vssd1 vccd1 vccd1 _2007_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2909_ _2355_/B hold740/X _2910_/S vssd1 vssd1 vccd1 vccd1 _2909_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2782__S hold38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2022__S _2055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2692__S _2697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2008__A1 _2036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold78_A hold78/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2625_ _2358_/B hold626/X _2633_/S vssd1 vssd1 vccd1 vccd1 _2625_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2556_ _2574_/A _2556_/B vssd1 vssd1 vccd1 vccd1 _2556_/X sky130_fd_sc_hd__and2_1
X_2487_ _1908_/D _2486_/X _2479_/X vssd1 vssd1 vccd1 vccd1 _2487_/X sky130_fd_sc_hd__a21o_2
XANTENNA__2867__S _2870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3108_ _3112_/A vssd1 vssd1 vccd1 vccd1 _3108_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_37_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3574_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3039_ _3049_/A vssd1 vssd1 vccd1 vccd1 _3039_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2777__S _2779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput25 hold1/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__clkbuf_1
Xinput36 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _1607_/A sky130_fd_sc_hd__clkbuf_2
Xinput14 input14/A vssd1 vssd1 vccd1 vccd1 _1612_/A sky130_fd_sc_hd__clkbuf_1
Xhold809 _1902_/Y vssd1 vssd1 vccd1 vccd1 hold809/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2410_ hold63/A hold20/A vssd1 vssd1 vccd1 vccd1 _2410_/X sky130_fd_sc_hd__and2_1
X_3390_ _3408_/CLK _3390_/D vssd1 vssd1 vccd1 vccd1 _3390_/Q sky130_fd_sc_hd__dfxtp_1
X_2341_ _3567_/Q _3566_/Q _3565_/Q _3564_/Q vssd1 vssd1 vccd1 vccd1 _2341_/X sky130_fd_sc_hd__or4_1
XFILLER_0_20_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2272_ _2272_/A _2278_/B vssd1 vssd1 vccd1 vccd1 _2275_/B sky130_fd_sc_hd__and2_1
XFILLER_0_79_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1987_ _2315_/A1 _1982_/X _1986_/X vssd1 vssd1 vccd1 vccd1 _1988_/A sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout122_A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2608_ _2103_/Y hold766/X _2612_/S vssd1 vssd1 vccd1 vccd1 _2608_/X sky130_fd_sc_hd__mux2_1
X_3588_ _3607_/CLK _3588_/D _3079_/Y vssd1 vssd1 vccd1 vccd1 _3588_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2539_ _3627_/Q hold11/A _2536_/X _2538_/X _2559_/B vssd1 vssd1 vccd1 vccd1 _2539_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_65_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_84_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2890_ _2058_/X hold676/X _2890_/S vssd1 vssd1 vccd1 vccd1 _2890_/X sky130_fd_sc_hd__mux2_1
X_1910_ _2162_/B hold470/X _1935_/A vssd1 vssd1 vccd1 vccd1 _1911_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_56_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1841_ _1877_/B vssd1 vssd1 vccd1 vccd1 _1841_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_60_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1772_ _1886_/A _1772_/B _1742_/B _1818_/A vssd1 vssd1 vccd1 vccd1 _1795_/B sky130_fd_sc_hd__or4bb_1
Xhold617 _2910_/X vssd1 vssd1 vccd1 vccd1 _3438_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold606 _3177_/Q vssd1 vssd1 vccd1 vccd1 hold606/X sky130_fd_sc_hd__dlygate4sd3_1
X_3511_ _3614_/CLK _3511_/D _3005_/Y vssd1 vssd1 vccd1 vccd1 _3511_/Q sky130_fd_sc_hd__dfrtp_1
X_3442_ _3589_/CLK _3442_/D _2936_/Y vssd1 vssd1 vccd1 vccd1 _3442_/Q sky130_fd_sc_hd__dfrtp_1
Xhold639 _2887_/X vssd1 vssd1 vccd1 vccd1 _3417_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 _3162_/Q vssd1 vssd1 vccd1 vccd1 hold628/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ _3413_/CLK _3373_/D vssd1 vssd1 vccd1 vccd1 _3373_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _2324_/A _2324_/B vssd1 vssd1 vccd1 vccd1 _2325_/C sky130_fd_sc_hd__xnor2_2
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2255_ _3466_/Q _2249_/A _3462_/Q vssd1 vssd1 vccd1 vccd1 _2255_/X sky130_fd_sc_hd__mux2_1
X_2186_ _2211_/A _2227_/A vssd1 vssd1 vccd1 vccd1 _2186_/X sky130_fd_sc_hd__or2_1
XANTENNA__2545__S1 _1943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2870__A1 _2356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2880__S _2880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2481__S0 _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2689__A1 _2801_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_52_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3408_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3650__A _3655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2040_ _2225_/A _2040_/B vssd1 vssd1 vccd1 vccd1 _2040_/X sky130_fd_sc_hd__and2b_1
X_2942_ _3122_/A vssd1 vssd1 vccd1 vccd1 _2942_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2873_ _2098_/S hold692/X _2880_/S vssd1 vssd1 vccd1 vccd1 _2873_/X sky130_fd_sc_hd__mux2_1
X_1824_ _1824_/A _1824_/B vssd1 vssd1 vccd1 vccd1 _3548_/D sky130_fd_sc_hd__nor2_1
X_1755_ _1811_/S _1755_/B _1769_/B vssd1 vssd1 vccd1 vccd1 _1755_/X sky130_fd_sc_hd__or3_1
XANTENNA__2463__S0 _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold403 _3261_/Q vssd1 vssd1 vccd1 vccd1 hold403/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 _2587_/X vssd1 vssd1 vccd1 vccd1 _3136_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 _2809_/X vssd1 vssd1 vccd1 vccd1 _3333_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 _3225_/Q vssd1 vssd1 vccd1 vccd1 hold425/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold458 _2214_/X vssd1 vssd1 vccd1 vccd1 _3481_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 _3491_/Q vssd1 vssd1 vccd1 vccd1 _1922_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold447 _3135_/Q vssd1 vssd1 vccd1 vccd1 hold447/X sky130_fd_sc_hd__dlygate4sd3_1
X_1686_ hold147/X _2399_/A hold65/X vssd1 vssd1 vccd1 vccd1 _1686_/X sky130_fd_sc_hd__mux2_1
X_3425_ _3431_/CLK _3425_/D vssd1 vssd1 vccd1 vccd1 _3425_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3356_ _3413_/CLK _3356_/D vssd1 vssd1 vccd1 vccd1 _3356_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _3484_/CLK _3287_/D vssd1 vssd1 vccd1 vccd1 _3287_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2875__S _2880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2307_ _1564_/Y _2064_/A _2041_/Y vssd1 vssd1 vccd1 vccd1 _2309_/A sky130_fd_sc_hd__a21oi_1
X_2238_ _2238_/A _2238_/B vssd1 vssd1 vccd1 vccd1 _2238_/Y sky130_fd_sc_hd__nor2_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2518__S1 _2532_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2169_ _2708_/A hold36/X _2168_/Y _2177_/A vssd1 vssd1 vccd1 vccd1 _2169_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold970 _1762_/X vssd1 vssd1 vccd1 vccd1 _3559_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 _3350_/Q vssd1 vssd1 vccd1 vccd1 _2146_/A sky130_fd_sc_hd__clkbuf_2
Xhold992 _1802_/Y vssd1 vssd1 vccd1 vccd1 hold992/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2785__S hold38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2598__A0 _2360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3210_ _3504_/CLK _3210_/D vssd1 vssd1 vccd1 vccd1 _3210_/Q sky130_fd_sc_hd__dfxtp_1
X_3141_ _3434_/CLK _3141_/D vssd1 vssd1 vccd1 vccd1 _3141_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2695__S _2697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3072_ _3097_/A vssd1 vssd1 vccd1 vccd1 _3072_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_82_45 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2825__A1 _2104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2023_ _2023_/A _2144_/C vssd1 vssd1 vccd1 vccd1 _2023_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2925_ _3127_/A vssd1 vssd1 vccd1 vccd1 _2925_/Y sky130_fd_sc_hd__inv_2
X_2856_ _2104_/B hold738/X _2860_/S vssd1 vssd1 vccd1 vccd1 _2856_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1807_ _1808_/A _3149_/Q vssd1 vssd1 vccd1 vccd1 _1886_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_60_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold200 _3287_/Q vssd1 vssd1 vccd1 vccd1 hold200/X sky130_fd_sc_hd__dlygate4sd3_1
X_2787_ _2807_/A1 hold368/X hold38/X vssd1 vssd1 vccd1 vccd1 _2787_/X sky130_fd_sc_hd__mux2_1
Xhold211 _2661_/X vssd1 vssd1 vccd1 vccd1 _3202_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2761__A0 _2801_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1738_ _1739_/A _1739_/B _1739_/C _1739_/D vssd1 vssd1 vccd1 vccd1 _1950_/C sky130_fd_sc_hd__nor4_1
Xhold233 _3314_/Q vssd1 vssd1 vccd1 vccd1 hold233/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _2804_/X vssd1 vssd1 vccd1 vccd1 _3328_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 _3137_/Q vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 _2791_/X vssd1 vssd1 vccd1 vccd1 _3316_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold255 _3253_/Q vssd1 vssd1 vccd1 vccd1 hold255/X sky130_fd_sc_hd__dlygate4sd3_1
X_1669_ _2401_/A _3606_/Q _1672_/S vssd1 vssd1 vccd1 vccd1 _1669_/X sky130_fd_sc_hd__mux2_1
Xhold277 _2735_/X vssd1 vssd1 vccd1 vccd1 _3266_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 _3289_/Q vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3408_ _3408_/CLK _3408_/D vssd1 vssd1 vccd1 vccd1 _3408_/Q sky130_fd_sc_hd__dfxtp_1
Xhold299 _3224_/Q vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _3408_/CLK _3339_/D vssd1 vssd1 vccd1 vccd1 _3339_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2816__A1 _2360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2427__S0 _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2807__A1 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2710_ _2801_/A1 hold220/X _2718_/S vssd1 vssd1 vccd1 vccd1 _2710_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2641_ _2357_/B hold666/X _2643_/S vssd1 vssd1 vccd1 vccd1 _2641_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2743__A0 _2803_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2572_ _2572_/A hold11/A _2572_/C _2572_/D vssd1 vssd1 vccd1 vccd1 _2574_/C sky130_fd_sc_hd__and4_1
XANTENNA__1607__B _1607_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1623__A hold92/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3124_ _3124_/A vssd1 vssd1 vccd1 vccd1 _3124_/Y sky130_fd_sc_hd__inv_2
X_3055_ _3057_/A vssd1 vssd1 vccd1 vccd1 _3055_/Y sky130_fd_sc_hd__inv_2
X_2006_ _3248_/Q _3320_/Q _3311_/Q _3302_/Q _2221_/B _2219_/A vssd1 vssd1 vccd1 vccd1
+ _2006_/X sky130_fd_sc_hd__mux4_1
X_2908_ _2357_/B hold592/X _2910_/S vssd1 vssd1 vccd1 vccd1 _2908_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2839_ _2356_/B hold732/X _2839_/S vssd1 vssd1 vccd1 vccd1 _2839_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1708__A _1767_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2725__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3330_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_output46_A _2571_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2624_ _3520_/Q _3519_/Q _2871_/C _2891_/B vssd1 vssd1 vccd1 vccd1 _2633_/S sky130_fd_sc_hd__or4b_4
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2716__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2555_ _2572_/C _2553_/X _2554_/X _2510_/B _3449_/Q vssd1 vssd1 vccd1 vccd1 _2556_/B
+ sky130_fd_sc_hd__a32o_1
X_2486_ _2485_/X _2482_/X _3518_/Q vssd1 vssd1 vccd1 vccd1 _2486_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2883__S _2890_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3107_ _3112_/A vssd1 vssd1 vccd1 vccd1 _3107_/Y sky130_fd_sc_hd__inv_2
X_3038_ _3067_/A vssd1 vssd1 vccd1 vccd1 _3038_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2707__A0 _2406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2793__S _2799_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput26 hold55/X vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__buf_1
XFILLER_0_64_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput37 wbs_we_i vssd1 vssd1 vccd1 vccd1 _1608_/A sky130_fd_sc_hd__clkbuf_2
Xinput15 hold17/X vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__2033__S _2055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3653__A _3655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2340_ _3563_/Q _3562_/Q _3561_/Q _3560_/Q vssd1 vssd1 vccd1 vccd1 _2340_/X sky130_fd_sc_hd__or4_1
XFILLER_0_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2271_ _2271_/A _2271_/B _2281_/B vssd1 vssd1 vccd1 vccd1 _2278_/B sky130_fd_sc_hd__and3_1
XANTENNA__1921__A1 _1918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2477__A2 hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1986_ _2315_/A1 _1986_/B vssd1 vssd1 vccd1 vccd1 _1986_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout115_A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2607_ _2105_/A hold712/X _2612_/S vssd1 vssd1 vccd1 vccd1 _2607_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2878__S _2880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3587_ _3600_/CLK _3587_/D _3078_/Y vssd1 vssd1 vccd1 vccd1 _3587_/Q sky130_fd_sc_hd__dfrtp_1
X_2538_ hold68/A _2438_/B _2572_/C _2537_/X vssd1 vssd1 vccd1 vccd1 _2538_/X sky130_fd_sc_hd__o211a_1
X_2469_ _2468_/X _2465_/X _3518_/Q vssd1 vssd1 vccd1 vccd1 _2469_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2788__S hold38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1840_ _1840_/A _3525_/Q _3524_/Q _3523_/Q vssd1 vssd1 vccd1 vccd1 _1877_/B sky130_fd_sc_hd__and4_2
XANTENNA__3648__A _3655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3510_ _3614_/CLK _3510_/D _3004_/Y vssd1 vssd1 vccd1 vccd1 _3510_/Q sky130_fd_sc_hd__dfrtp_1
X_1771_ _1771_/A _1771_/B _3552_/Q vssd1 vssd1 vccd1 vccd1 _1798_/C sky130_fd_sc_hd__and3_1
XFILLER_0_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold618 _3168_/Q vssd1 vssd1 vccd1 vccd1 hold618/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold607 _2630_/X vssd1 vssd1 vccd1 vccd1 _3177_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3441_ _3589_/CLK _3441_/D _2935_/Y vssd1 vssd1 vccd1 vccd1 _3441_/Q sky130_fd_sc_hd__dfrtp_1
Xhold629 _2612_/X vssd1 vssd1 vccd1 vccd1 _3162_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _3579_/CLK _3372_/D vssd1 vssd1 vccd1 vccd1 _3372_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _2323_/A _2323_/B vssd1 vssd1 vccd1 vccd1 _2324_/B sky130_fd_sc_hd__xnor2_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2254_ _3467_/Q hold852/X _3462_/Q vssd1 vssd1 vccd1 vccd1 _2254_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_18_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2185_ _2211_/A _2182_/Y _2184_/X vssd1 vssd1 vccd1 vccd1 _2227_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1969_ hold196/X hold222/X hold192/X hold208/X _2045_/S0 _2045_/S1 vssd1 vssd1 vccd1
+ vccd1 _1969_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_50_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2481__S1 _1943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1992__S0 _2045_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2356__B _2356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_21_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3633_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2074__B1 _2355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1983__S0 _2221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2301__A1 hold75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2941_ _3032_/A vssd1 vssd1 vccd1 vccd1 _2941_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2872_ _2358_/B hold758/X _2880_/S vssd1 vssd1 vccd1 vccd1 _2872_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_37_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1823_ _1810_/Y _1818_/B _1818_/A vssd1 vssd1 vccd1 vccd1 _1823_/Y sky130_fd_sc_hd__a21oi_1
X_1754_ hold979/X _2387_/C _1753_/X vssd1 vssd1 vccd1 vccd1 _1754_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_13_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2463__S1 _1943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold404 _2728_/X vssd1 vssd1 vccd1 vccd1 _3261_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold415 _3331_/Q vssd1 vssd1 vccd1 vccd1 hold415/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 _2687_/X vssd1 vssd1 vccd1 vccd1 _3225_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1685_ hold323/X _2400_/A hold65/X vssd1 vssd1 vccd1 vccd1 _3594_/D sky130_fd_sc_hd__mux2_1
X_3424_ _3424_/CLK _3424_/D vssd1 vssd1 vccd1 vccd1 _3424_/Q sky130_fd_sc_hd__dfxtp_1
Xhold437 _3243_/Q vssd1 vssd1 vccd1 vccd1 hold437/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 _2586_/X vssd1 vssd1 vccd1 vccd1 _3135_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 _3478_/Q vssd1 vssd1 vccd1 vccd1 hold459/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3355_ _3413_/CLK _3355_/D vssd1 vssd1 vccd1 vccd1 _3355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _3605_/CLK _3286_/D vssd1 vssd1 vccd1 vccd1 _3286_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ _1564_/Y _2065_/B _1999_/A vssd1 vssd1 vccd1 vccd1 _2310_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__2540__A1 _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2237_ _2259_/B _2240_/A vssd1 vssd1 vccd1 vccd1 _2237_/Y sky130_fd_sc_hd__nor2_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2168_ hold36/X _2225_/B vssd1 vssd1 vccd1 vccd1 _2168_/Y sky130_fd_sc_hd__nand2_1
X_2099_ _2099_/A _2099_/B vssd1 vssd1 vccd1 vccd1 _2111_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold971 _3566_/Q vssd1 vssd1 vccd1 vccd1 hold971/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold982 _2386_/X vssd1 vssd1 vccd1 vccd1 _3350_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold960 _1770_/X vssd1 vssd1 vccd1 vccd1 _3556_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 _1804_/Y vssd1 vssd1 vccd1 vccd1 _3553_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3140_ _3434_/CLK _3140_/D vssd1 vssd1 vccd1 vccd1 _3140_/Q sky130_fd_sc_hd__dfxtp_1
X_3071_ _3097_/A vssd1 vssd1 vccd1 vccd1 _3071_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_82_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2022_ _2023_/A _2021_/X _2055_/S vssd1 vssd1 vccd1 vccd1 _2022_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1612__C _1624_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2589__A1 _2406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2924_ _3127_/A vssd1 vssd1 vccd1 vccd1 _2924_/Y sky130_fd_sc_hd__inv_2
X_2855_ _2105_/A hold754/X _2860_/S vssd1 vssd1 vccd1 vccd1 _2855_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1806_ _1806_/A1 _1798_/D hold834/X vssd1 vssd1 vccd1 vccd1 _1806_/Y sky130_fd_sc_hd__a21oi_1
Xhold201 _2758_/X vssd1 vssd1 vccd1 vccd1 _3287_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2786_ _2806_/A1 hold263/X hold38/X vssd1 vssd1 vccd1 vccd1 _2786_/X sky130_fd_sc_hd__mux2_1
X_1737_ _1581_/Y _3452_/Q hold83/X _1585_/Y _1730_/X vssd1 vssd1 vccd1 vccd1 _1739_/D
+ sky130_fd_sc_hd__a221o_1
Xhold234 _2788_/X vssd1 vssd1 vccd1 vccd1 _3314_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 _3206_/Q vssd1 vssd1 vccd1 vccd1 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 _2588_/X vssd1 vssd1 vccd1 vccd1 _3137_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _3280_/Q vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 _3294_/Q vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 _2720_/X vssd1 vssd1 vccd1 vccd1 _3253_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 _3325_/Q vssd1 vssd1 vccd1 vccd1 hold278/X sky130_fd_sc_hd__dlygate4sd3_1
X_1668_ hold98/A _1668_/B vssd1 vssd1 vccd1 vccd1 _1668_/Y sky130_fd_sc_hd__nand2_1
Xhold289 _2761_/X vssd1 vssd1 vccd1 vccd1 _3289_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3407_ _3434_/CLK _3407_/D vssd1 vssd1 vccd1 vccd1 _3407_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2886__S _2890_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3338_ _3434_/CLK _3338_/D vssd1 vssd1 vccd1 vccd1 _3338_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1599_ _2146_/A vssd1 vssd1 vccd1 vccd1 _1599_/Y sky130_fd_sc_hd__inv_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3269_ _3484_/CLK _3269_/D vssd1 vssd1 vccd1 vccd1 _3269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2427__S1 _1943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2752__A1 _2802_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2796__S _2799_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold790 _3507_/Q vssd1 vssd1 vccd1 vccd1 hold790/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2268__B1 _2270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2036__S _2036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2640_ _2360_/B hold572/X _2643_/S vssd1 vssd1 vccd1 vccd1 _2640_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2571_ _3454_/Q hold35/A hold20/A vssd1 vssd1 vccd1 vccd1 _2571_/X sky130_fd_sc_hd__and3_2
XFILLER_0_77_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1623__B input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3123_ _3124_/A vssd1 vssd1 vccd1 vccd1 _3123_/Y sky130_fd_sc_hd__inv_2
X_3054_ _3054_/A vssd1 vssd1 vccd1 vccd1 _3054_/Y sky130_fd_sc_hd__inv_2
X_2005_ _3293_/Q _3284_/Q _3275_/Q _3266_/Q _2221_/B _2219_/A vssd1 vssd1 vccd1 vccd1
+ _2005_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2907_ _2360_/B hold576/X _2910_/S vssd1 vssd1 vccd1 vccd1 _2907_/X sky130_fd_sc_hd__mux2_1
X_2838_ _2355_/B hold522/X _2839_/S vssd1 vssd1 vccd1 vccd1 _2838_/X sky130_fd_sc_hd__mux2_1
X_2769_ hold30/X _2769_/A1 _2769_/S vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__mux2_1
XFILLER_0_13_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2734__A1 _2804_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2498__B1 _2492_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output39_A _3439_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2661__A0 _2804_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2623_ _2356_/B hold670/X _2623_/S vssd1 vssd1 vccd1 vccd1 _2623_/X sky130_fd_sc_hd__mux2_1
X_2554_ _3589_/Q _2558_/B _2438_/B _3601_/Q vssd1 vssd1 vccd1 vccd1 _2554_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_2_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2485_ _2484_/X _2483_/X _3517_/Q vssd1 vssd1 vccd1 vccd1 _2485_/X sky130_fd_sc_hd__mux2_1
X_3106_ _3129_/A vssd1 vssd1 vccd1 vccd1 _3106_/Y sky130_fd_sc_hd__inv_2
X_3037_ _3067_/A vssd1 vssd1 vccd1 vccd1 _3037_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2652__A0 _2357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_46_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3521_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2359__B _2360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2643__A0 _2356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput27 input27/A vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_1
Xinput16 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 _1624_/B sky130_fd_sc_hd__buf_2
XFILLER_0_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2270_ _2270_/A _2270_/B _2270_/C vssd1 vssd1 vccd1 vccd1 _2281_/B sky130_fd_sc_hd__and3_1
XANTENNA__2269__B _2270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1685__A1 _2400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_2_0__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1985_ _1984_/X _1983_/X _2036_/S vssd1 vssd1 vccd1 vccd1 _1986_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_7_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3655_ _3655_/A vssd1 vssd1 vccd1 vccd1 _3655_/X sky130_fd_sc_hd__buf_1
XFILLER_0_70_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2606_ _2109_/B hold714/X _2612_/S vssd1 vssd1 vccd1 vccd1 _2606_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout108_A hold120/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3586_ _3589_/CLK _3586_/D _3077_/Y vssd1 vssd1 vccd1 vccd1 _3586_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2537_ _3587_/Q _2558_/B _2558_/C _3381_/Q vssd1 vssd1 vccd1 vccd1 _2537_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2468_ _2467_/X _2466_/X _2546_/S vssd1 vssd1 vccd1 vccd1 _2468_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2894__S _2900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2399_ _2399_/A hold98/X hold95/X vssd1 vssd1 vccd1 vccd1 _3581_/D sky130_fd_sc_hd__and3_1
XANTENNA__2873__A0 _2098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2625__A0 _2358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2616__A0 _2098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2044__S _2055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1770_ hold959/X _2387_/C _1769_/X vssd1 vssd1 vccd1 vccd1 _1770_/X sky130_fd_sc_hd__o21a_1
Xhold608 _3432_/Q vssd1 vssd1 vccd1 vccd1 hold608/X sky130_fd_sc_hd__dlygate4sd3_1
X_3440_ _3589_/CLK _3440_/D _2934_/Y vssd1 vssd1 vccd1 vccd1 _3440_/Q sky130_fd_sc_hd__dfrtp_1
Xhold619 _2620_/X vssd1 vssd1 vccd1 vccd1 _3168_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3371_ _3431_/CLK _3371_/D vssd1 vssd1 vccd1 vccd1 _3371_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2322_ _2322_/A _2322_/B vssd1 vssd1 vccd1 vccd1 _2323_/B sky130_fd_sc_hd__xnor2_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2253_ hold858/X _3467_/Q _3462_/Q vssd1 vssd1 vccd1 vccd1 _2253_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1912__A _2546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2855__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2184_ _2184_/A _2211_/A hold36/X _2198_/B vssd1 vssd1 vccd1 vccd1 _2184_/X sky130_fd_sc_hd__or4_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__2607__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1968_ hold780/X _1967_/Y _2055_/S vssd1 vssd1 vccd1 vccd1 _1968_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2889__S _2890_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1899_ _1904_/A _2613_/B vssd1 vssd1 vccd1 vccd1 _1905_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_43_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3638_ _3638_/CLK _3638_/D _3129_/Y vssd1 vssd1 vccd1 vccd1 _3638_/Q sky130_fd_sc_hd__dfrtp_1
X_3569_ _3573_/CLK _3569_/D _3063_/Y vssd1 vssd1 vccd1 vccd1 _3569_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1992__S1 _2045_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1649__A1 hold70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1968__S _2055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2799__S _2799_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1983__S1 _2195_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2837__A0 _2357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2940_ _3032_/A vssd1 vssd1 vccd1 vccd1 _2940_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_84_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2871_ _3520_/Q _3519_/Q _2871_/C _2901_/B vssd1 vssd1 vccd1 vccd1 _2880_/S sky130_fd_sc_hd__or4b_4
XFILLER_0_57_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1822_ _1742_/B _1824_/A _1821_/Y _1814_/B vssd1 vssd1 vccd1 vccd1 _3549_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_4_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1753_ _1811_/S _1753_/B _1769_/B vssd1 vssd1 vccd1 vccd1 _1753_/X sky130_fd_sc_hd__or3_1
XFILLER_0_4_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold416 _2807_/X vssd1 vssd1 vccd1 vccd1 _3331_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 _3205_/Q vssd1 vssd1 vccd1 vccd1 hold427/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold405 _3134_/Q vssd1 vssd1 vccd1 vccd1 hold405/X sky130_fd_sc_hd__dlygate4sd3_1
X_1684_ hold128/X _2401_/A hold65/X vssd1 vssd1 vccd1 vccd1 _3595_/D sky130_fd_sc_hd__mux2_1
X_3423_ _3579_/CLK _3423_/D vssd1 vssd1 vccd1 vccd1 _3423_/Q sky130_fd_sc_hd__dfxtp_1
Xhold438 _2707_/X vssd1 vssd1 vccd1 vccd1 _3243_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 _3212_/Q vssd1 vssd1 vccd1 vccd1 hold449/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _3413_/CLK _3354_/D vssd1 vssd1 vccd1 vccd1 _3354_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ hold338/X _2576_/A hold22/X vssd1 vssd1 vccd1 vccd1 _3440_/D sky130_fd_sc_hd__mux2_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ _3321_/CLK _3285_/D vssd1 vssd1 vccd1 vccd1 _3285_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2236_ _2259_/A _2238_/A _2230_/B vssd1 vssd1 vccd1 vccd1 _2236_/X sky130_fd_sc_hd__o21ba_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2167_ _2708_/A _2171_/A vssd1 vssd1 vccd1 vccd1 _2225_/B sky130_fd_sc_hd__xnor2_1
X_2098_ _2358_/B _2095_/Y _2098_/S vssd1 vssd1 vccd1 vccd1 _2099_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_61_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold972 _1748_/X vssd1 vssd1 vccd1 vccd1 _3566_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 _3561_/Q vssd1 vssd1 vccd1 vccd1 _1755_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold950 _1820_/X vssd1 vssd1 vccd1 vccd1 _3550_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 _3536_/Q vssd1 vssd1 vccd1 vccd1 _1859_/A sky130_fd_sc_hd__buf_1
Xhold994 _3148_/Q vssd1 vssd1 vccd1 vccd1 hold994/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3070_ _3101_/A vssd1 vssd1 vccd1 vccd1 _3070_/Y sky130_fd_sc_hd__inv_2
X_2021_ _3505_/Q _2144_/C _2020_/X vssd1 vssd1 vccd1 vccd1 _2021_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_82_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2923_ _3049_/A vssd1 vssd1 vccd1 vccd1 _2923_/Y sky130_fd_sc_hd__inv_2
X_2854_ _2109_/B hold632/X _2860_/S vssd1 vssd1 vccd1 vccd1 _2854_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1805_ _1772_/B _1798_/D _3552_/Q vssd1 vssd1 vccd1 vccd1 _1805_/Y sky130_fd_sc_hd__a21oi_1
X_2785_ _2805_/A1 hold301/X hold38/X vssd1 vssd1 vccd1 vccd1 _2785_/X sky130_fd_sc_hd__mux2_1
Xhold202 _3269_/Q vssd1 vssd1 vccd1 vccd1 hold202/X sky130_fd_sc_hd__dlygate4sd3_1
X_1736_ _1736_/A _1736_/B _1736_/C _1736_/D vssd1 vssd1 vccd1 vccd1 _2381_/B sky130_fd_sc_hd__or4_4
Xhold224 _3262_/Q vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 _2665_/X vssd1 vssd1 vccd1 vccd1 _3206_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 _3490_/Q vssd1 vssd1 vccd1 vccd1 _2708_/A sky130_fd_sc_hd__buf_2
Xhold246 _2751_/X vssd1 vssd1 vccd1 vccd1 _3280_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 _2766_/X vssd1 vssd1 vccd1 vccd1 _3294_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1667_ _1667_/A _2413_/A vssd1 vssd1 vccd1 vccd1 _2437_/A sky130_fd_sc_hd__nor2_2
Xhold257 _3489_/Q vssd1 vssd1 vccd1 vccd1 _2729_/B sky130_fd_sc_hd__buf_2
X_3406_ _3433_/CLK _3406_/D vssd1 vssd1 vccd1 vccd1 _3406_/Q sky130_fd_sc_hd__dfxtp_1
X_1598_ _1957_/B vssd1 vssd1 vccd1 vccd1 _1598_/Y sky130_fd_sc_hd__inv_2
Xhold279 _2801_/X vssd1 vssd1 vccd1 vccd1 _3325_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3337_ _3433_/CLK _3337_/D vssd1 vssd1 vccd1 vccd1 _3337_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2513__A2 hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _3321_/CLK _3268_/D vssd1 vssd1 vccd1 vccd1 _3268_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2187__B _2219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3199_ _3330_/CLK _3199_/D vssd1 vssd1 vccd1 vccd1 _3199_/Q sky130_fd_sc_hd__dfxtp_1
X_2219_ _2219_/A _2219_/B vssd1 vssd1 vccd1 vccd1 _2223_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold791 _1990_/X vssd1 vssd1 vccd1 vccd1 _3507_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold780 _3509_/Q vssd1 vssd1 vccd1 vccd1 hold780/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2268__A1 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2570_ _2574_/A _2570_/B vssd1 vssd1 vccd1 vccd1 _2570_/X sky130_fd_sc_hd__and2_1
X_3122_ _3122_/A vssd1 vssd1 vccd1 vccd1 _3122_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1623__C _1623_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3053_ _3054_/A vssd1 vssd1 vccd1 vccd1 _3053_/Y sky130_fd_sc_hd__inv_2
X_2004_ _3221_/Q _3212_/Q _3203_/Q _3329_/Q _2045_/S0 _2045_/S1 vssd1 vssd1 vccd1
+ vccd1 _2004_/X sky130_fd_sc_hd__mux4_1
X_2906_ _2104_/B hold654/X _2910_/S vssd1 vssd1 vccd1 vccd1 _2906_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2837_ _2357_/B hold558/X _2839_/S vssd1 vssd1 vccd1 vccd1 _2837_/X sky130_fd_sc_hd__mux2_1
X_2768_ _2808_/A1 hold204/X _2769_/S vssd1 vssd1 vccd1 vccd1 _2768_/X sky130_fd_sc_hd__mux2_1
X_1719_ _1853_/A _3454_/Q vssd1 vssd1 vccd1 vccd1 _1719_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__2897__S _2900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2699_ _2801_/A1 hold407/X _2707_/S vssd1 vssd1 vccd1 vccd1 _2699_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2498__A1 _1908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2670__A1 _2803_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2571__A _3454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2622_ _2355_/B hold662/X _2623_/S vssd1 vssd1 vccd1 vccd1 _2622_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2553_ hold67/A hold11/A _2558_/C _3383_/Q _2559_/B vssd1 vssd1 vccd1 vccd1 _2553_/X
+ sky130_fd_sc_hd__o221a_1
X_2484_ _3175_/Q _3424_/Q _3415_/Q _3157_/Q _1918_/B _1912_/B vssd1 vssd1 vccd1 vccd1
+ _2484_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2024__S0 _2045_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3105_ _3110_/A vssd1 vssd1 vccd1 vccd1 _3105_/Y sky130_fd_sc_hd__inv_2
X_3036_ _3067_/A vssd1 vssd1 vccd1 vccd1 _3036_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1915__B1 _2546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3594_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2015__S0 _2045_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput17 hold61/X vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__clkbuf_2
Xinput28 input28/A vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_1
XANTENNA__1719__B _3454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2006__S0 _2221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1613__C_N _1623_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2505__S _3518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1984_ _3250_/Q _3322_/Q _3313_/Q _3304_/Q _2221_/B _2219_/A vssd1 vssd1 vccd1 vccd1
+ _1984_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2493__S0 _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3654_ _3655_/A vssd1 vssd1 vccd1 vccd1 _3654_/X sky130_fd_sc_hd__buf_1
XFILLER_0_70_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2605_ _2098_/S hold612/X _2612_/S vssd1 vssd1 vccd1 vccd1 _2605_/X sky130_fd_sc_hd__mux2_1
X_3585_ _3600_/CLK _3585_/D _3076_/Y vssd1 vssd1 vccd1 vccd1 _3585_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2536_ _3618_/Q _1643_/Y hold11/A vssd1 vssd1 vccd1 vccd1 _2536_/X sky130_fd_sc_hd__a21bo_1
X_2467_ _3174_/Q _3423_/Q _3414_/Q _3156_/Q _2532_/S0 _1912_/B vssd1 vssd1 vccd1 vccd1
+ _2467_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2398_ _2576_/A hold98/X hold95/X vssd1 vssd1 vccd1 vccd1 _3580_/D sky130_fd_sc_hd__and3_1
XFILLER_0_3_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3019_ _3057_/A vssd1 vssd1 vccd1 vccd1 _3019_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2484__S0 _1918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1555__A _1767_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2864__A1 _2109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold609 _2904_/X vssd1 vssd1 vccd1 vccd1 _3432_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3370_ _3424_/CLK _3370_/D vssd1 vssd1 vccd1 vccd1 _3370_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2321_ _2321_/A _2321_/B vssd1 vssd1 vccd1 vccd1 _2322_/B sky130_fd_sc_hd__xnor2_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2252_ hold862/X hold858/X _3462_/Q vssd1 vssd1 vccd1 vccd1 _2252_/X sky130_fd_sc_hd__mux2_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1912__B _1912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2183_ hold36/X _2198_/B vssd1 vssd1 vccd1 vccd1 _2183_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2466__S0 _2532_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1967_ _2144_/C _1967_/B vssd1 vssd1 vccd1 vccd1 _1967_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout120_A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1898_ _1891_/A _2613_/B _1897_/Y _1924_/A vssd1 vssd1 vccd1 vccd1 _1898_/X sky130_fd_sc_hd__o211a_1
X_3637_ _3638_/CLK _3637_/D _3128_/Y vssd1 vssd1 vccd1 vccd1 _3637_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3568_ _3573_/CLK _3568_/D _3062_/Y vssd1 vssd1 vccd1 vccd1 _3568_/Q sky130_fd_sc_hd__dfrtp_1
X_2519_ _3178_/Q _3427_/Q _3418_/Q _3160_/Q _1918_/B _2532_/S1 vssd1 vssd1 vccd1 vccd1
+ _2519_/X sky130_fd_sc_hd__mux4_1
X_3499_ _3555_/CLK _3499_/D _2993_/Y vssd1 vssd1 vccd1 vccd1 _3499_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2074__A2 _2357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2782__A0 _2802_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3638_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2870_ hold494/X _2356_/B _2870_/S vssd1 vssd1 vccd1 vccd1 _2870_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2055__S _2055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1821_ _1742_/B _1818_/A _1810_/A vssd1 vssd1 vccd1 vccd1 _1821_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1752_ _1749_/B _2387_/C _1751_/X vssd1 vssd1 vccd1 vccd1 _1752_/X sky130_fd_sc_hd__o21a_1
Xhold406 _2585_/X vssd1 vssd1 vccd1 vccd1 _3134_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 _3232_/Q vssd1 vssd1 vccd1 vccd1 hold417/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1683_ hold85/X hold75/X hold65/X vssd1 vssd1 vccd1 vccd1 _3596_/D sky130_fd_sc_hd__mux2_1
X_3422_ _3579_/CLK _3422_/D vssd1 vssd1 vccd1 vccd1 _3422_/Q sky130_fd_sc_hd__dfxtp_1
Xhold428 _2664_/X vssd1 vssd1 vccd1 vccd1 _3205_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 _3204_/Q vssd1 vssd1 vccd1 vccd1 hold439/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _3431_/CLK _3353_/D vssd1 vssd1 vccd1 vccd1 _3353_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _3319_/CLK _3284_/D vssd1 vssd1 vccd1 vccd1 _3284_/Q sky130_fd_sc_hd__dfxtp_1
X_2304_ _1724_/B _2399_/A hold22/X vssd1 vssd1 vccd1 vccd1 _3441_/D sky130_fd_sc_hd__mux2_1
X_2235_ _2259_/B _2240_/A vssd1 vssd1 vccd1 vccd1 _2238_/A sky130_fd_sc_hd__and2_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2828__A1 _2355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2166_ _2729_/B _3488_/Q _2677_/B vssd1 vssd1 vccd1 vccd1 _2171_/A sky130_fd_sc_hd__and3_1
X_2097_ _2095_/A _2095_/B _2096_/Y vssd1 vssd1 vccd1 vccd1 _2097_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_75_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2999_ _3101_/A vssd1 vssd1 vccd1 vccd1 _2999_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_71_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2764__A0 _2804_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold940 _3349_/Q vssd1 vssd1 vccd1 vccd1 hold940/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 _1758_/X vssd1 vssd1 vccd1 vccd1 _3561_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold951 _3560_/Q vssd1 vssd1 vccd1 vccd1 _1757_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 _3151_/Q vssd1 vssd1 vccd1 vccd1 _1809_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold984 _1860_/X vssd1 vssd1 vccd1 vccd1 _3536_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 _3459_/Q vssd1 vssd1 vccd1 vccd1 _2271_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2819__A1 _2356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1979__S _2055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2383__B _2383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2020_ _2315_/A1 _2018_/X _2019_/X _2014_/X _2000_/S vssd1 vssd1 vccd1 vccd1 _2020_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_82_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2574__A _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2922_ _3127_/A vssd1 vssd1 vccd1 vccd1 _2922_/Y sky130_fd_sc_hd__inv_2
X_2853_ _2098_/S hold750/X _2860_/S vssd1 vssd1 vccd1 vccd1 _2853_/X sky130_fd_sc_hd__mux2_1
X_1804_ _1798_/D _1803_/X hold992/X vssd1 vssd1 vccd1 vccd1 _1804_/Y sky130_fd_sc_hd__a21oi_1
X_2784_ _2804_/A1 hold145/X hold38/X vssd1 vssd1 vccd1 vccd1 _2784_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2746__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1735_ _1736_/A _1736_/B _1736_/C _1736_/D vssd1 vssd1 vccd1 vccd1 _1950_/B sky130_fd_sc_hd__nor4_1
XFILLER_0_25_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold225 _2731_/X vssd1 vssd1 vccd1 vccd1 _3262_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 _2738_/X vssd1 vssd1 vccd1 vccd1 _3269_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold214 _3133_/Q vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 _3298_/Q vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__dlygate4sd3_1
X_1666_ _1666_/A _2421_/A vssd1 vssd1 vccd1 vccd1 _2418_/B sky130_fd_sc_hd__nand2_1
Xhold258 _2173_/X vssd1 vssd1 vccd1 vccd1 _3489_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 _2169_/X vssd1 vssd1 vccd1 vccd1 _3490_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 _3441_/Q vssd1 vssd1 vccd1 vccd1 _1724_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3405_ _3434_/CLK _3405_/D vssd1 vssd1 vccd1 vccd1 _3405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1597_ _2144_/C vssd1 vssd1 vccd1 vccd1 _2000_/S sky130_fd_sc_hd__inv_2
X_3336_ _3434_/CLK _3336_/D vssd1 vssd1 vccd1 vccd1 _3336_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _3321_/CLK _3267_/D vssd1 vssd1 vccd1 vccd1 _3267_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2187__C _2221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3198_ _3424_/CLK _3198_/D vssd1 vssd1 vccd1 vccd1 _3198_/Q sky130_fd_sc_hd__dfxtp_1
X_2218_ _3488_/Q _3487_/Q vssd1 vssd1 vccd1 vccd1 _2219_/B sky130_fd_sc_hd__xor2_1
X_2149_ _2146_/A _2381_/D _2146_/B vssd1 vssd1 vccd1 vccd1 _2157_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold770 _3190_/Q vssd1 vssd1 vccd1 vccd1 hold770/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 _1968_/X vssd1 vssd1 vccd1 vccd1 _3509_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 _3503_/Q vssd1 vssd1 vccd1 vccd1 hold792/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold929_A _3439_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2728__A0 _2406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3121_ _3124_/A vssd1 vssd1 vccd1 vccd1 _3121_/Y sky130_fd_sc_hd__inv_2
X_3052_ _3054_/A vssd1 vssd1 vccd1 vccd1 _3052_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_26_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2003_ _2036_/S _2003_/B vssd1 vssd1 vccd1 vccd1 _2003_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2905_ _2105_/A hold582/X _2910_/S vssd1 vssd1 vccd1 vccd1 _2905_/X sky130_fd_sc_hd__mux2_1
X_2836_ _2360_/B hold636/X _2839_/S vssd1 vssd1 vccd1 vccd1 _2836_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2195__A1 _2195_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2767_ _2807_/A1 hold330/X _2769_/S vssd1 vssd1 vccd1 vccd1 _2767_/X sky130_fd_sc_hd__mux2_1
X_1718_ hold83/A _1877_/A vssd1 vssd1 vccd1 vccd1 _1718_/X sky130_fd_sc_hd__and2b_1
X_2698_ _2719_/A hold37/X vssd1 vssd1 vccd1 vccd1 _2707_/S sky130_fd_sc_hd__or2_4
X_1649_ _3616_/Q hold70/X hold53/X vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__mux2_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2198__B _2198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ _3319_/CLK _3319_/D vssd1 vssd1 vccd1 vccd1 _3319_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2621_ _2357_/B hold554/X _2623_/S vssd1 vssd1 vccd1 vccd1 _2621_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2552_ _1908_/D _2547_/X _2549_/X _2551_/X vssd1 vssd1 vccd1 vccd1 _2552_/X sky130_fd_sc_hd__a211o_2
XFILLER_0_23_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2483_ _3374_/Q _3356_/Q _3365_/Q _3193_/Q _2532_/S0 _2532_/S1 vssd1 vssd1 vccd1
+ vccd1 _2483_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2024__S1 _2045_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3104_ _3112_/A vssd1 vssd1 vccd1 vccd1 _3104_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_37_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3035_ _3067_/A vssd1 vssd1 vccd1 vccd1 _3035_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2184__D _2198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2819_ hold584/X _2356_/B _2819_/S vssd1 vssd1 vccd1 vccd1 _2819_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2701__S _2707_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1915__A1 _1912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2015__S1 _2045_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput18 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 _1657_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_52_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput29 input29/A vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_1
XANTENNA__2611__S _2612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2006__S1 _2219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output44_A _2567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1983_ _3295_/Q _3286_/Q _3277_/Q _3268_/Q _2221_/B _2195_/A1 vssd1 vssd1 vccd1 vccd1
+ _1983_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2493__S1 _1943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3653_ _3655_/A vssd1 vssd1 vccd1 vccd1 _3653_/X sky130_fd_sc_hd__buf_1
XFILLER_0_70_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2604_ _2358_/B hold722/X _2612_/S vssd1 vssd1 vccd1 vccd1 _2604_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2521__S _3518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3584_ _3600_/CLK _3584_/D _3075_/Y vssd1 vssd1 vccd1 vccd1 _3584_/Q sky130_fd_sc_hd__dfrtp_1
X_2535_ hold73/A hold35/A hold20/A vssd1 vssd1 vccd1 vccd1 _2535_/X sky130_fd_sc_hd__and3_1
XFILLER_0_11_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2466_ _3373_/Q _3355_/Q _3364_/Q _3192_/Q _2532_/S0 _1912_/B vssd1 vssd1 vccd1 vccd1
+ _2466_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_48_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2397_ hold94/A hold63/A vssd1 vssd1 vccd1 vccd1 _2558_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_78_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3018_ _3054_/A vssd1 vssd1 vccd1 vccd1 _3018_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2484__S1 _1912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2606__S _2612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2552__A1 _1908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2320_ _1564_/Y _1785_/Y _2009_/X vssd1 vssd1 vccd1 vccd1 _2321_/B sky130_fd_sc_hd__a21oi_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2251_ _2248_/A _3469_/Q _3462_/Q vssd1 vssd1 vccd1 vccd1 _2251_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2304__A1 _2399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1912__C _1918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2182_ _2375_/B vssd1 vssd1 vccd1 vccd1 _2182_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_0_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3326_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1966_ _2315_/A1 _1961_/X _1965_/X vssd1 vssd1 vccd1 vccd1 _1967_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__2466__S1 _1912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2791__A1 _2801_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1897_ _2613_/B _1946_/B vssd1 vssd1 vccd1 vccd1 _1897_/Y sky130_fd_sc_hd__nand2_1
X_3636_ _3638_/CLK _3636_/D _3127_/Y vssd1 vssd1 vccd1 vccd1 _3636_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout113_A hold123/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3567_ _3567_/CLK _3567_/D _3061_/Y vssd1 vssd1 vccd1 vccd1 _3567_/Q sky130_fd_sc_hd__dfstp_1
X_2518_ _3377_/Q _3359_/Q _3368_/Q _3196_/Q _2532_/S0 _2532_/S1 vssd1 vssd1 vccd1
+ vccd1 _2518_/X sky130_fd_sc_hd__mux4_1
X_3498_ _3555_/CLK _3498_/D _2992_/Y vssd1 vssd1 vccd1 vccd1 _3498_/Q sky130_fd_sc_hd__dfrtp_1
X_2449_ _3372_/Q _3354_/Q _3363_/Q _3191_/Q _2532_/S0 _2532_/S1 vssd1 vssd1 vccd1
+ vccd1 _2449_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_66_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2950__A _3124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold7 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1820_ _1772_/B hold949/X _1815_/X vssd1 vssd1 vccd1 vccd1 _1820_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_44_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2773__A1 _2803_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1751_ _1811_/S _3563_/Q _1769_/B vssd1 vssd1 vccd1 vccd1 _1751_/X sky130_fd_sc_hd__or3_1
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold418 _2695_/X vssd1 vssd1 vccd1 vccd1 _3232_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold407 _3235_/Q vssd1 vssd1 vccd1 vccd1 hold407/X sky130_fd_sc_hd__dlygate4sd3_1
X_1682_ hold82/X hold70/X hold65/X vssd1 vssd1 vccd1 vccd1 _3597_/D sky130_fd_sc_hd__mux2_1
X_3421_ _3424_/CLK _3421_/D vssd1 vssd1 vccd1 vccd1 _3421_/Q sky130_fd_sc_hd__dfxtp_1
Xhold429 _3214_/Q vssd1 vssd1 vccd1 vccd1 hold429/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1959__S0 _2045_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3352_ _3550_/CLK _3352_/D _2927_/Y vssd1 vssd1 vccd1 vccd1 _3352_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ _1726_/B _2400_/A hold22/X vssd1 vssd1 vccd1 vccd1 _3442_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _3332_/CLK _3283_/D vssd1 vssd1 vccd1 vccd1 _3283_/Q sky130_fd_sc_hd__dfxtp_1
X_2234_ _2234_/A _2234_/B vssd1 vssd1 vccd1 vccd1 _2234_/X sky130_fd_sc_hd__and2_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2165_ hold35/X _2165_/B _2165_/C vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__and3_1
X_2096_ _2096_/A _2096_/B vssd1 vssd1 vccd1 vccd1 _2096_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_0_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2998_ _3101_/A vssd1 vssd1 vccd1 vccd1 _2998_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_9_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1949_ _3510_/Q _1948_/Y hold471/X vssd1 vssd1 vccd1 vccd1 _1949_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_71_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3619_ _3619_/CLK _3619_/D _3110_/Y vssd1 vssd1 vccd1 vccd1 _3619_/Q sky130_fd_sc_hd__dfrtp_1
Xhold930 _3494_/Q vssd1 vssd1 vccd1 vccd1 _2130_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 _3458_/Q vssd1 vssd1 vccd1 vccd1 _2271_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold952 _1760_/X vssd1 vssd1 vccd1 vccd1 _3560_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 _2371_/X vssd1 vssd1 vccd1 vccd1 hold941/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 _2278_/Y vssd1 vssd1 vccd1 vccd1 _3459_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 hold985/A vssd1 vssd1 vccd1 vccd1 _2157_/A sky130_fd_sc_hd__buf_1
Xhold974 _1794_/X vssd1 vssd1 vccd1 vccd1 _3150_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2755__A1 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2921_ _3127_/A vssd1 vssd1 vccd1 vccd1 _2921_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2852_ _2358_/B hold682/X _2860_/S vssd1 vssd1 vccd1 vccd1 _2852_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2783_ _2803_/A1 hold327/X hold38/X vssd1 vssd1 vccd1 vccd1 _2783_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1918__B _1918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1803_ _1771_/B _3552_/Q _1600_/Y vssd1 vssd1 vccd1 vccd1 _1803_/X sky130_fd_sc_hd__a21o_1
X_1734_ _1879_/A hold173/X _1718_/X _1721_/X _1724_/X vssd1 vssd1 vccd1 vccd1 _1736_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_79_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold204 _3296_/Q vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 _3271_/Q vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 _2584_/X vssd1 vssd1 vccd1 vccd1 _3133_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold259 _3307_/Q vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__dlygate4sd3_1
X_3404_ _3431_/CLK _3404_/D vssd1 vssd1 vccd1 vccd1 _3404_/Q sky130_fd_sc_hd__dfxtp_1
Xhold237 _3220_/Q vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
X_1665_ _1574_/A _2576_/A _1665_/S vssd1 vssd1 vccd1 vccd1 _3607_/D sky130_fd_sc_hd__mux2_1
Xhold248 _3607_/Q vssd1 vssd1 vccd1 vccd1 _1574_/A sky130_fd_sc_hd__dlygate4sd3_1
X_1596_ _3345_/Q vssd1 vssd1 vccd1 vccd1 _1596_/Y sky130_fd_sc_hd__inv_2
X_3335_ _3434_/CLK _3335_/D vssd1 vssd1 vccd1 vccd1 _3335_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ _3320_/CLK _3266_/D vssd1 vssd1 vccd1 vccd1 _3266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2217_ _2211_/Y _2211_/B _2217_/S vssd1 vssd1 vccd1 vccd1 _2217_/X sky130_fd_sc_hd__mux2_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3197_ _3516_/CLK _3197_/D vssd1 vssd1 vccd1 vccd1 _3197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2682__A0 _2804_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2148_ _2375_/A _2148_/B vssd1 vssd1 vccd1 vccd1 _2158_/S sky130_fd_sc_hd__nand2_1
X_2079_ _2070_/A _2078_/X _2076_/X vssd1 vssd1 vccd1 vccd1 _2079_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_48_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1788__A2 _2064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2704__S _2707_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2737__A1 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold771 _2646_/X vssd1 vssd1 vccd1 vccd1 _3190_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold760 _3167_/Q vssd1 vssd1 vccd1 vccd1 hold760/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout93_A _2195_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold782 _3502_/Q vssd1 vssd1 vccd1 vccd1 _2053_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold793 _2033_/X vssd1 vssd1 vccd1 vccd1 _3503_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3120_ _3122_/A vssd1 vssd1 vccd1 vccd1 _3120_/Y sky130_fd_sc_hd__inv_2
X_3051_ _3054_/A vssd1 vssd1 vccd1 vccd1 _3051_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2664__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2002_ _3257_/Q _3134_/Q _3239_/Q _3230_/Q _2045_/S0 _2045_/S1 vssd1 vssd1 vccd1
+ vccd1 _2003_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_18_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2904_ _2109_/B hold608/X _2910_/S vssd1 vssd1 vccd1 vccd1 _2904_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2835_ _2104_/B hold764/X _2839_/S vssd1 vssd1 vccd1 vccd1 _2835_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2766_ _2806_/A1 hold267/X _2769_/S vssd1 vssd1 vccd1 vccd1 _2766_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1717_ _1848_/A _1717_/B vssd1 vssd1 vccd1 vccd1 _1717_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2697_ hold445/X _2406_/A _2697_/S vssd1 vssd1 vccd1 vccd1 _2697_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1648_ hold90/X hold87/X hold53/X vssd1 vssd1 vccd1 vccd1 _3617_/D sky130_fd_sc_hd__mux2_1
X_3318_ _3318_/CLK _3318_/D vssd1 vssd1 vccd1 vccd1 _3318_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1579_ _3540_/Q vssd1 vssd1 vccd1 vccd1 _1579_/Y sky130_fd_sc_hd__inv_2
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3249_ _3321_/CLK _3249_/D vssd1 vssd1 vccd1 vccd1 _3249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2502__S0 _1918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold590 _3379_/Q vssd1 vssd1 vccd1 vccd1 hold590/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2609__S _2612_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2646__A0 _2358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1621__A1 _2399_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2620_ _2360_/B hold618/X _2623_/S vssd1 vssd1 vccd1 vccd1 _2620_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2551_ _3619_/Q _1643_/Y _2510_/B _3448_/Q _2550_/Y vssd1 vssd1 vccd1 vccd1 _2551_/X
+ sky130_fd_sc_hd__a221o_1
X_2482_ _2481_/X _2480_/X _2546_/S vssd1 vssd1 vccd1 vccd1 _2482_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2885__A0 _2101_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3103_ _3110_/A vssd1 vssd1 vccd1 vccd1 _3103_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2637__A0 _2109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3034_ _3069_/A vssd1 vssd1 vccd1 vccd1 _3034_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_73_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2818_ hold674/X _2355_/B _2819_/S vssd1 vssd1 vccd1 vccd1 _2818_/X sky130_fd_sc_hd__mux2_1
X_2749_ _2406_/A hold349/X _2749_/S vssd1 vssd1 vccd1 vccd1 _2749_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2573__C1 _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1915__A2 _1918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2876__A0 _2104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1679__A1 _2406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2429__S _2546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2628__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2953__A _3124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3533_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_64_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput19 hold97/X vssd1 vssd1 vccd1 vccd1 _1607_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2619__A0 _2104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1982_ _1980_/X _1981_/X _2036_/S vssd1 vssd1 vccd1 vccd1 _1982_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3652_ _3655_/A vssd1 vssd1 vccd1 vccd1 _3652_/X sky130_fd_sc_hd__buf_1
X_2603_ _2901_/A _2891_/B vssd1 vssd1 vccd1 vccd1 _2612_/S sky130_fd_sc_hd__nand2_4
X_3583_ _3610_/CLK _3583_/D _3074_/Y vssd1 vssd1 vccd1 vccd1 _3583_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2534_ _2533_/X _2530_/X _3518_/Q vssd1 vssd1 vccd1 vccd1 _2534_/X sky130_fd_sc_hd__mux2_1
X_2465_ _2464_/X _2463_/X _2546_/S vssd1 vssd1 vccd1 vccd1 _2465_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2858__A0 _2357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2396_ hold94/X hold63/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__and2_1
X_3017_ _3032_/A vssd1 vssd1 vccd1 vccd1 _3017_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2712__S _2718_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1995__S1 _2219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2849__A0 _2356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3019__A _3057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ _3466_/Q _2247_/X _2249_/X hold846/X vssd1 vssd1 vccd1 vccd1 _2250_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_20_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2181_ _2144_/A _2180_/X _2372_/S vssd1 vssd1 vccd1 vccd1 _2198_/B sky130_fd_sc_hd__o21bai_4
XFILLER_0_79_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1965_ _2315_/A1 _1965_/B vssd1 vssd1 vccd1 vccd1 _1965_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1896_ _1896_/A _1896_/B vssd1 vssd1 vccd1 vccd1 _1946_/B sky130_fd_sc_hd__or2_1
XFILLER_0_43_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3635_ _3635_/CLK _3635_/D _3126_/Y vssd1 vssd1 vccd1 vccd1 _3635_/Q sky130_fd_sc_hd__dfrtp_1
X_3566_ _3567_/CLK _3566_/D _3060_/Y vssd1 vssd1 vccd1 vccd1 _3566_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout106_A hold117/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2517_ _2516_/X _2515_/X _2546_/S vssd1 vssd1 vccd1 vccd1 _2517_/X sky130_fd_sc_hd__mux2_1
X_3497_ _3555_/CLK _3497_/D _2991_/Y vssd1 vssd1 vccd1 vccd1 _3497_/Q sky130_fd_sc_hd__dfrtp_1
X_2448_ _2447_/X _2446_/X _2546_/S vssd1 vssd1 vccd1 vccd1 _2448_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2379_ _2379_/A _2379_/B _2379_/C vssd1 vssd1 vccd1 vccd1 _2379_/X sky130_fd_sc_hd__and3_1
XANTENNA__2707__S _2707_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2298__A1 hold45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__buf_1
XFILLER_0_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2470__A1 _1908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1750_ _1747_/B _2387_/C _1749_/X vssd1 vssd1 vccd1 vccd1 _1750_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_80_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1681_ _3598_/Q hold87/X hold65/X vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__mux2_1
XFILLER_0_20_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold408 _2699_/X vssd1 vssd1 vccd1 vccd1 _3235_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3420_ _3424_/CLK _3420_/D vssd1 vssd1 vccd1 vccd1 _3420_/Q sky130_fd_sc_hd__dfxtp_1
Xhold419 _3591_/Q vssd1 vssd1 vccd1 vccd1 _2211_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1959__S1 _2045_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2525__A2 hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3351_ _3550_/CLK _3351_/D _2926_/Y vssd1 vssd1 vccd1 vccd1 _3351_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2302_ hold173/X _2401_/A hold22/X vssd1 vssd1 vccd1 vccd1 _3443_/D sky130_fd_sc_hd__mux2_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _3318_/CLK _3282_/D vssd1 vssd1 vccd1 vccd1 _3282_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2233_ _2232_/A _2230_/B _2230_/A vssd1 vssd1 vccd1 vccd1 _2233_/X sky130_fd_sc_hd__a21o_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2164_ _3478_/Q _3577_/Q hold98/A vssd1 vssd1 vccd1 vccd1 _2165_/C sky130_fd_sc_hd__and3b_1
X_2095_ _2095_/A _2095_/B vssd1 vssd1 vccd1 vccd1 _2095_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2997_ _3101_/A vssd1 vssd1 vccd1 vccd1 _2997_/Y sky130_fd_sc_hd__inv_2
X_1948_ _3518_/Q _1893_/B _1932_/B _1945_/Y _1947_/Y vssd1 vssd1 vccd1 vccd1 _1948_/Y
+ sky130_fd_sc_hd__a2111oi_1
X_1879_ _1879_/A _1879_/B vssd1 vssd1 vccd1 vccd1 _1879_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold920 _3513_/Q vssd1 vssd1 vccd1 vccd1 _1929_/A sky130_fd_sc_hd__dlygate4sd3_1
X_3618_ _3627_/CLK hold54/X _3109_/Y vssd1 vssd1 vccd1 vccd1 _3618_/Q sky130_fd_sc_hd__dfrtp_1
Xhold931 _2153_/X vssd1 vssd1 vccd1 vccd1 hold931/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 _2280_/X vssd1 vssd1 vccd1 vccd1 _3458_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 _3558_/Q vssd1 vssd1 vccd1 vccd1 _1761_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold942 _2372_/X vssd1 vssd1 vccd1 vccd1 _3348_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 hold997/A vssd1 vssd1 vccd1 vccd1 _2119_/B sky130_fd_sc_hd__buf_1
X_3549_ _3559_/CLK _3549_/D _3043_/Y vssd1 vssd1 vccd1 vccd1 _3549_/Q sky130_fd_sc_hd__dfrtp_1
Xhold986 _2381_/X vssd1 vssd1 vccd1 vccd1 hold986/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 _3551_/Q vssd1 vssd1 vccd1 vccd1 _1886_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2010__B _2144_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2900__S _2900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2140__B1 _2000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2691__A1 _2803_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2920_ _3097_/A vssd1 vssd1 vccd1 vccd1 _2920_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2851_ _2881_/B _2901_/B vssd1 vssd1 vccd1 vccd1 _2860_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_38_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2782_ _2802_/A1 hold129/X hold38/X vssd1 vssd1 vccd1 vccd1 _2782_/X sky130_fd_sc_hd__mux2_1
X_1802_ _3552_/Q _1798_/D _1771_/B vssd1 vssd1 vccd1 vccd1 _1802_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1733_ _1879_/A hold173/X _1717_/Y _1720_/Y _1722_/Y vssd1 vssd1 vccd1 vccd1 _1736_/C
+ sky130_fd_sc_hd__o2111ai_2
Xhold205 _2768_/X vssd1 vssd1 vccd1 vccd1 _3296_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 _3487_/Q vssd1 vssd1 vccd1 vccd1 _2677_/B sky130_fd_sc_hd__clkbuf_2
Xhold227 _2741_/X vssd1 vssd1 vccd1 vccd1 _3271_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 _3249_/Q vssd1 vssd1 vccd1 vccd1 hold249/X sky130_fd_sc_hd__dlygate4sd3_1
X_3403_ _3438_/CLK _3403_/D vssd1 vssd1 vccd1 vccd1 _3403_/Q sky130_fd_sc_hd__dfxtp_1
Xhold238 _2682_/X vssd1 vssd1 vccd1 vccd1 _3220_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1664_ _1573_/A _2399_/A _1665_/S vssd1 vssd1 vccd1 vccd1 _3608_/D sky130_fd_sc_hd__mux2_1
X_1595_ _3346_/Q vssd1 vssd1 vccd1 vccd1 _1595_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3334_ _3432_/CLK _3334_/D vssd1 vssd1 vccd1 vccd1 _3334_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _3332_/CLK _3265_/D vssd1 vssd1 vccd1 vccd1 _3265_/Q sky130_fd_sc_hd__dfxtp_1
X_2216_ _2204_/B _2211_/Y _2215_/X _2211_/B _2202_/A vssd1 vssd1 vccd1 vccd1 _2216_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3196_ _3619_/CLK _3196_/D vssd1 vssd1 vccd1 vccd1 _3196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2147_ _1957_/B _2379_/B _2155_/C vssd1 vssd1 vccd1 vccd1 _2148_/B sky130_fd_sc_hd__mux2_1
X_2078_ _2068_/Y _2077_/Y _2092_/A vssd1 vssd1 vccd1 vccd1 _2078_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2434__A1 _1908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2720__S _2728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_49_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3432_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold750 _3386_/Q vssd1 vssd1 vccd1 vccd1 hold750/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 _3164_/Q vssd1 vssd1 vccd1 vccd1 hold772/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold761 _2619_/X vssd1 vssd1 vccd1 vccd1 _3167_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2045__S0 _2045_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout86_A _2532_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold794 _3506_/Q vssd1 vssd1 vccd1 vccd1 _2010_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 _2044_/X vssd1 vssd1 vccd1 vccd1 _3502_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2673__A1 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2630__S _2633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3050_ _3054_/A vssd1 vssd1 vccd1 vccd1 _3050_/Y sky130_fd_sc_hd__inv_2
X_2001_ _2010_/A _2000_/X _2055_/S vssd1 vssd1 vccd1 vccd1 _2001_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2903_ _2098_/S hold716/X _2910_/S vssd1 vssd1 vccd1 vccd1 _2903_/X sky130_fd_sc_hd__mux2_1
X_2834_ _2101_/Y hold600/X _2839_/S vssd1 vssd1 vccd1 vccd1 _2834_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2765_ _2805_/A1 hold351/X _2769_/S vssd1 vssd1 vccd1 vccd1 _2765_/X sky130_fd_sc_hd__mux2_1
X_1716_ _3534_/Q _1716_/B vssd1 vssd1 vccd1 vccd1 _1716_/Y sky130_fd_sc_hd__nand2b_1
X_2696_ hold208/X _2808_/A1 _2697_/S vssd1 vssd1 vccd1 vccd1 _2696_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2027__S0 _2221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1647_ _3618_/Q hold45/X hold53/X vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__mux2_1
XFILLER_0_41_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1578_ _3603_/Q vssd1 vssd1 vccd1 vccd1 _1578_/Y sky130_fd_sc_hd__inv_2
X_3317_ _3319_/CLK _3317_/D vssd1 vssd1 vccd1 vccd1 _3317_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _3320_/CLK _3248_/D vssd1 vssd1 vccd1 vccd1 _3248_/Q sky130_fd_sc_hd__dfxtp_1
X_3179_ _3579_/CLK _3179_/D vssd1 vssd1 vccd1 vccd1 _3179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2715__S _2718_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2502__S1 _1912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold580 _3197_/Q vssd1 vssd1 vccd1 vccd1 hold580/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 _2849_/X vssd1 vssd1 vccd1 vccd1 _3379_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1590__A _2221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2625__S _2633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2550_ _2550_/A hold11/A vssd1 vssd1 vccd1 vccd1 _2550_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_23_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2481_ _3184_/Q _3337_/Q _3166_/Q _3142_/Q _1944_/B _1943_/A vssd1 vssd1 vccd1 vccd1
+ _2481_/X sky130_fd_sc_hd__mux4_1
X_3102_ _3112_/A vssd1 vssd1 vccd1 vccd1 _3102_/Y sky130_fd_sc_hd__inv_2
X_3033_ _3069_/A vssd1 vssd1 vccd1 vccd1 _3033_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2496__S0 _1918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2817_ hold492/X _2357_/B _2819_/S vssd1 vssd1 vccd1 vccd1 _2817_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2748_ _2808_/A1 hold188/X _2749_/S vssd1 vssd1 vccd1 vccd1 _2748_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2679_ _2801_/A1 hold261/X _2687_/S vssd1 vssd1 vccd1 vccd1 _2679_/X sky130_fd_sc_hd__mux2_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2867__A1 _2360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1751__C _1769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1981_ hold411/X hold429/X hold427/X hold415/X _2045_/S0 _2045_/S1 vssd1 vssd1 vccd1
+ vccd1 _1981_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_55_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3651_ _3655_/A vssd1 vssd1 vccd1 vccd1 _3651_/X sky130_fd_sc_hd__buf_1
X_3582_ _3590_/CLK _3582_/D _3073_/Y vssd1 vssd1 vccd1 vccd1 _3582_/Q sky130_fd_sc_hd__dfrtp_1
X_2602_ _3522_/Q _3521_/Q vssd1 vssd1 vccd1 vccd1 _2891_/B sky130_fd_sc_hd__nor2_4
X_2533_ _2532_/X _2531_/X _3517_/Q vssd1 vssd1 vccd1 vccd1 _2533_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2464_ _3183_/Q _3336_/Q _3165_/Q _3141_/Q _1944_/B _1943_/A vssd1 vssd1 vccd1 vccd1
+ _2464_/X sky130_fd_sc_hd__mux4_1
X_2395_ _2395_/A _2395_/B _2395_/C vssd1 vssd1 vccd1 vccd1 _2395_/X sky130_fd_sc_hd__or3_2
X_3016_ _3110_/A vssd1 vssd1 vccd1 vccd1 _3016_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_80_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout120 input2/X vssd1 vssd1 vccd1 vccd1 _3112_/A sky130_fd_sc_hd__buf_8
XFILLER_0_69_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2785__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2180_ _2490_/A _3348_/Q vssd1 vssd1 vccd1 vccd1 _2180_/X sky130_fd_sc_hd__and2_1
X_1964_ _1963_/X _1962_/X _2222_/A vssd1 vssd1 vccd1 vccd1 _1965_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1895_ _1902_/A _3519_/Q _1891_/A vssd1 vssd1 vccd1 vccd1 _1896_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3634_ _3638_/CLK _3634_/D _3125_/Y vssd1 vssd1 vccd1 vccd1 _3634_/Q sky130_fd_sc_hd__dfrtp_1
X_3565_ _3567_/CLK _3565_/D _3059_/Y vssd1 vssd1 vccd1 vccd1 _3565_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2516_ _3187_/Q _3340_/Q _3169_/Q _3145_/Q _2532_/S0 _2532_/S1 vssd1 vssd1 vccd1
+ vccd1 _2516_/X sky130_fd_sc_hd__mux4_1
X_3496_ _3550_/CLK _3496_/D _2990_/Y vssd1 vssd1 vccd1 vccd1 _3496_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2447_ _3182_/Q _3335_/Q _3164_/Q _3140_/Q _1944_/B _1943_/A vssd1 vssd1 vccd1 vccd1
+ _2447_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_75_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2700__A0 _2802_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2378_ _2378_/A1 _2370_/A _2377_/X _2144_/D _2372_/S vssd1 vssd1 vccd1 vccd1 _2378_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2767__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2723__S _2728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__buf_1
XFILLER_0_71_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2633__S _2633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold409 _3138_/Q vssd1 vssd1 vccd1 vccd1 hold409/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1680_ hold68/X hold45/X hold65/X vssd1 vssd1 vccd1 vccd1 _3599_/D sky130_fd_sc_hd__mux2_1
X_3350_ _3635_/CLK _3350_/D _2925_/Y vssd1 vssd1 vccd1 vccd1 _3350_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2301_ hold83/X hold75/X hold22/X vssd1 vssd1 vccd1 vccd1 _3444_/D sky130_fd_sc_hd__mux2_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _3322_/CLK _3281_/D vssd1 vssd1 vccd1 vccd1 _3281_/Q sky130_fd_sc_hd__dfxtp_1
X_2232_ _2232_/A _3476_/Q vssd1 vssd1 vccd1 vccd1 _2259_/D sky130_fd_sc_hd__nor2_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2163_ _1922_/A _1929_/B _2162_/X _1935_/A vssd1 vssd1 vccd1 vccd1 _2163_/X sky130_fd_sc_hd__a211o_1
X_2094_ _2064_/B _2091_/X _2093_/X _2067_/B vssd1 vssd1 vccd1 vccd1 _2095_/B sky130_fd_sc_hd__a211oi_1
XANTENNA__2109__A _2360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2543__S _2546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2749__A0 _2406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2996_ _3101_/A vssd1 vssd1 vccd1 vccd1 _2996_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_56_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1947_ _3518_/Q _1893_/B _1946_/X vssd1 vssd1 vccd1 vccd1 _1947_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1878_ _1837_/A _1842_/Y _1877_/X _1877_/A _1836_/A vssd1 vssd1 vccd1 vccd1 _1878_/X
+ sky130_fd_sc_hd__a32o_1
Xhold921 _3567_/Q vssd1 vssd1 vccd1 vccd1 hold921/X sky130_fd_sc_hd__dlygate4sd3_1
X_3617_ _3622_/CLK _3617_/D _3108_/Y vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold910 _3153_/Q vssd1 vssd1 vccd1 vccd1 _1808_/D sky130_fd_sc_hd__buf_1
Xhold954 _1764_/X vssd1 vssd1 vccd1 vccd1 _3558_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3548_ _3559_/CLK _3548_/D _3042_/Y vssd1 vssd1 vccd1 vccd1 _3548_/Q sky130_fd_sc_hd__dfrtp_1
Xhold932 _2154_/X vssd1 vssd1 vccd1 vccd1 _3494_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 hold943/A vssd1 vssd1 vccd1 vccd1 _1957_/A sky130_fd_sc_hd__buf_1
Xhold998 _3532_/Q vssd1 vssd1 vccd1 vccd1 _1848_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold965 _3525_/Q vssd1 vssd1 vccd1 vccd1 _1839_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold987 _2382_/Y vssd1 vssd1 vccd1 vccd1 _3349_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 _1817_/X vssd1 vssd1 vccd1 vccd1 _3551_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3479_ _3605_/CLK _3479_/D _2973_/Y vssd1 vssd1 vccd1 vccd1 _3479_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__1659__A_N hold62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2718__S _2718_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2628__S _2633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2443__A2 hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2850_ _3522_/Q _3521_/Q vssd1 vssd1 vccd1 vccd1 _2901_/B sky130_fd_sc_hd__and2_2
XFILLER_0_5_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1801_ _1801_/A _1801_/B vssd1 vssd1 vccd1 vccd1 _1801_/X sky130_fd_sc_hd__and2_1
X_2781_ _2801_/A1 hold259/X hold38/X vssd1 vssd1 vccd1 vccd1 _2781_/X sky130_fd_sc_hd__mux2_1
X_1732_ _1580_/Y _3455_/Q _1709_/X _1710_/X _1712_/X vssd1 vssd1 vccd1 vccd1 _1736_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold206 _3229_/Q vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
X_1663_ _1572_/A _2400_/A _1665_/S vssd1 vssd1 vccd1 vccd1 _3609_/D sky130_fd_sc_hd__mux2_1
Xhold217 _2179_/X vssd1 vssd1 vccd1 vccd1 _3487_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 _3305_/Q vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
X_3402_ _3438_/CLK _3402_/D vssd1 vssd1 vccd1 vccd1 _3402_/Q sky130_fd_sc_hd__dfxtp_1
Xhold228 _3635_/Q vssd1 vssd1 vccd1 vccd1 _1950_/A sky130_fd_sc_hd__buf_1
X_1594_ _3458_/Q vssd1 vssd1 vccd1 vccd1 _1594_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2903__A0 _2098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _3333_/CLK _3333_/D vssd1 vssd1 vccd1 vccd1 _3333_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _3318_/CLK _3264_/D vssd1 vssd1 vccd1 vccd1 _3264_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2215_ _3479_/Q _2215_/B vssd1 vssd1 vccd1 vccd1 _2215_/X sky130_fd_sc_hd__or2_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _3516_/CLK _3195_/D vssd1 vssd1 vccd1 vccd1 _3195_/Q sky130_fd_sc_hd__dfxtp_1
X_2146_ _2146_/A _2146_/B vssd1 vssd1 vccd1 vccd1 _2155_/C sky130_fd_sc_hd__or2_1
X_2077_ _3544_/Q _2084_/B vssd1 vssd1 vccd1 vccd1 _2077_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2979_ _3097_/A vssd1 vssd1 vccd1 vccd1 _2979_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold751 _2853_/X vssd1 vssd1 vccd1 vccd1 _3386_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 _2616_/X vssd1 vssd1 vccd1 vccd1 _3164_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 _3165_/Q vssd1 vssd1 vccd1 vccd1 hold762/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold740 _3437_/Q vssd1 vssd1 vccd1 vccd1 hold740/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2045__S1 _2045_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold795 _2001_/X vssd1 vssd1 vccd1 vccd1 _3506_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 _3504_/Q vssd1 vssd1 vccd1 vccd1 _2023_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2448__S _2546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3607_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2000_ hold790/X _1999_/Y _2000_/S vssd1 vssd1 vccd1 vccd1 _2000_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2902_ _2358_/B hold724/X _2910_/S vssd1 vssd1 vccd1 vccd1 _2902_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2833_ _2109_/B hold644/X _2839_/S vssd1 vssd1 vccd1 vccd1 _2833_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2821__S _2829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2764_ _2804_/A1 hold155/X _2769_/S vssd1 vssd1 vccd1 vccd1 _2764_/X sky130_fd_sc_hd__mux2_1
X_1715_ _3451_/Q _1850_/A vssd1 vssd1 vccd1 vccd1 _1715_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2695_ hold417/X _2807_/A1 _2697_/S vssd1 vssd1 vccd1 vccd1 _2695_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2027__S1 _2219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1646_ hold396/X _2406_/A hold53/X vssd1 vssd1 vccd1 vccd1 _3619_/D sky130_fd_sc_hd__mux2_1
X_1577_ _3604_/Q vssd1 vssd1 vccd1 vccd1 _1577_/Y sky130_fd_sc_hd__inv_2
X_3316_ _3318_/CLK _3316_/D vssd1 vssd1 vccd1 vccd1 _3316_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ _3319_/CLK _3247_/D vssd1 vssd1 vccd1 vccd1 _3247_/Q sky130_fd_sc_hd__dfxtp_1
X_3178_ _3575_/CLK _3178_/D vssd1 vssd1 vccd1 vccd1 _3178_/Q sky130_fd_sc_hd__dfxtp_1
X_2129_ _2129_/A _2157_/A vssd1 vssd1 vccd1 vccd1 _2155_/B sky130_fd_sc_hd__or2_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold570 _3337_/Q vssd1 vssd1 vccd1 vccd1 hold570/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 _2653_/X vssd1 vssd1 vccd1 vccd1 _3197_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 _3436_/Q vssd1 vssd1 vccd1 vccd1 hold592/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1749__C _1769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2582__A1 _2802_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2480_ _3406_/Q _3397_/Q _3388_/Q _3433_/Q _1944_/B _1943_/A vssd1 vssd1 vccd1 vccd1
+ _2480_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3101_ _3101_/A vssd1 vssd1 vccd1 vccd1 _3101_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_37_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3032_ _3032_/A vssd1 vssd1 vccd1 vccd1 _3032_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2098__A0 _2358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2496__S1 _1912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2816_ hold544/X _2360_/B _2819_/S vssd1 vssd1 vccd1 vccd1 _2816_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1956__A _2144_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout129_A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2747_ _2807_/A1 hold370/X _2749_/S vssd1 vssd1 vccd1 vccd1 _2747_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2678_ _2800_/B _2760_/A vssd1 vssd1 vccd1 vccd1 _2687_/S sky130_fd_sc_hd__or2_4
X_1629_ hold27/X hold25/X hold12/X vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__mux2_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2726__S _2728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1630__S hold12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2025__A_N _2036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3555_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1827__A0 _2383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1980_ hold401/X hold435/X hold421/X hold417/X _2045_/S0 _2045_/S1 vssd1 vssd1 vccd1
+ vccd1 _1980_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_28_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3650_ _3655_/A vssd1 vssd1 vccd1 vccd1 _3650_/X sky130_fd_sc_hd__buf_1
XFILLER_0_70_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2601_ _2356_/B hold668/X _2601_/S vssd1 vssd1 vccd1 vccd1 _2601_/X sky130_fd_sc_hd__mux2_1
X_3581_ _3607_/CLK _3581_/D _3072_/Y vssd1 vssd1 vccd1 vccd1 _3581_/Q sky130_fd_sc_hd__dfrtp_1
X_2532_ _3179_/Q _3428_/Q _3419_/Q _3161_/Q _2532_/S0 _2532_/S1 vssd1 vssd1 vccd1
+ vccd1 _2532_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_23_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2463_ _3405_/Q _3396_/Q _3387_/Q _3432_/Q _1944_/B _1943_/A vssd1 vssd1 vccd1 vccd1
+ _2463_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_11_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2394_ _3601_/Q _3383_/Q _3345_/Q _3594_/Q _2392_/X vssd1 vssd1 vccd1 vccd1 _2395_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2400__A _2400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2546__S _2546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3015_ _3110_/A vssd1 vssd1 vccd1 vccd1 _3015_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_80_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2794__A1 _2804_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout121 input2/X vssd1 vssd1 vccd1 vccd1 _3090_/A sky130_fd_sc_hd__buf_8
Xfanout110 hold126/X vssd1 vssd1 vccd1 vccd1 _2802_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output42_A _2561_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1963_ hold357/X hold47/X _3315_/Q hold40/X _2049_/S0 _2219_/A vssd1 vssd1 vccd1
+ vccd1 _1963_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_28_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2776__A1 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1894_ _1892_/A _2613_/B _1893_/Y _1924_/A vssd1 vssd1 vccd1 vccd1 _1894_/X sky130_fd_sc_hd__o211a_1
X_3633_ _3633_/CLK hold28/X _3124_/Y vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfstp_1
XANTENNA__2114__B _2383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3564_ _3567_/CLK _3564_/D _3058_/Y vssd1 vssd1 vccd1 vccd1 _3564_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2515_ _3409_/Q _3400_/Q _3391_/Q _3436_/Q _1944_/B _1943_/A vssd1 vssd1 vccd1 vccd1
+ _2515_/X sky130_fd_sc_hd__mux4_1
X_3495_ _3635_/CLK _3495_/D _2989_/Y vssd1 vssd1 vccd1 vccd1 _3495_/Q sky130_fd_sc_hd__dfrtp_1
X_2446_ _3404_/Q _3395_/Q _3386_/Q _3431_/Q _1944_/B _1943_/A vssd1 vssd1 vccd1 vccd1
+ _2446_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2377_ _2379_/B _2379_/C _2377_/C vssd1 vssd1 vccd1 vccd1 _2377_/X sky130_fd_sc_hd__and3_1
XFILLER_0_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2975__A _3124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2758__A1 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1757__C _1769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3280_ _3321_/CLK _3280_/D vssd1 vssd1 vccd1 vccd1 _3280_/Q sky130_fd_sc_hd__dfxtp_1
X_2300_ hold84/X hold70/X hold22/X vssd1 vssd1 vccd1 vccd1 _3445_/D sky130_fd_sc_hd__mux2_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ _2232_/A _2234_/A vssd1 vssd1 vccd1 vccd1 _2231_/Y sky130_fd_sc_hd__xnor2_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2162_ _2871_/C _2162_/B _2162_/C vssd1 vssd1 vccd1 vccd1 _2162_/X sky130_fd_sc_hd__and3_1
X_2093_ _2092_/A _1579_/Y _2064_/A _2092_/Y vssd1 vssd1 vccd1 vccd1 _2093_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2541__S0 _1918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2109__B _2109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2824__S _2829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2995_ _3129_/A vssd1 vssd1 vccd1 vccd1 _2995_/Y sky130_fd_sc_hd__inv_2
X_1946_ _2546_/S _1946_/B vssd1 vssd1 vccd1 vccd1 _1946_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1877_ _1877_/A _1877_/B vssd1 vssd1 vccd1 vccd1 _1877_/X sky130_fd_sc_hd__or2_1
Xhold922 _1746_/X vssd1 vssd1 vccd1 vccd1 _3567_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold900 _3573_/Q vssd1 vssd1 vccd1 vccd1 _1698_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout111_A hold126/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3616_ _3627_/CLK hold71/X _3107_/Y vssd1 vssd1 vccd1 vccd1 _3616_/Q sky130_fd_sc_hd__dfrtp_1
Xhold911 _2376_/X vssd1 vssd1 vccd1 vccd1 _3153_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 _3565_/Q vssd1 vssd1 vccd1 vccd1 _1747_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 _3564_/Q vssd1 vssd1 vccd1 vccd1 _1749_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3547_ _3571_/CLK _3547_/D _3041_/Y vssd1 vssd1 vccd1 vccd1 _3547_/Q sky130_fd_sc_hd__dfrtp_1
Xhold933 _3496_/Q vssd1 vssd1 vccd1 vccd1 _2139_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold988 _3476_/Q vssd1 vssd1 vccd1 vccd1 _2230_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 _1882_/X vssd1 vssd1 vccd1 vccd1 _3525_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 _3548_/Q vssd1 vssd1 vccd1 vccd1 _1818_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold999 _1868_/X vssd1 vssd1 vccd1 vccd1 _3532_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3478_ _3590_/CLK _3478_/D _2972_/Y vssd1 vssd1 vccd1 vccd1 _3478_/Q sky130_fd_sc_hd__dfrtp_1
X_2429_ _2428_/X _2427_/X _2546_/S vssd1 vssd1 vccd1 vccd1 _2429_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2685__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2532__S0 _2532_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1651__A1 _2401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1800_ _1771_/B _3552_/Q _1798_/D _1771_/A vssd1 vssd1 vccd1 vccd1 _1800_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2780_ hold37/X _2790_/B vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__or2_1
X_1731_ _1584_/Y hold89/X hold338/X _1885_/S _1714_/X vssd1 vssd1 vccd1 vccd1 _1736_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2600__A0 _2355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold207 _2692_/X vssd1 vssd1 vccd1 vccd1 _3229_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1662_ _3610_/Q _2401_/A _1665_/S vssd1 vssd1 vccd1 vccd1 _1662_/X sky130_fd_sc_hd__mux2_1
Xhold218 _3251_/Q vssd1 vssd1 vccd1 vccd1 hold218/X sky130_fd_sc_hd__dlygate4sd3_1
X_3401_ _3521_/CLK _3401_/D vssd1 vssd1 vccd1 vccd1 _3401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold229 _1621_/X vssd1 vssd1 vccd1 vccd1 _3635_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1593_ _3459_/Q vssd1 vssd1 vccd1 vccd1 _1593_/Y sky130_fd_sc_hd__inv_2
X_3332_ _3332_/CLK _3332_/D vssd1 vssd1 vccd1 vccd1 _3332_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _3319_/CLK _3263_/D vssd1 vssd1 vccd1 vccd1 _3263_/Q sky130_fd_sc_hd__dfxtp_1
X_2214_ _2210_/B _2211_/Y _2213_/X _2211_/B _2205_/A vssd1 vssd1 vccd1 vccd1 _2214_/X
+ sky130_fd_sc_hd__a32o_1
X_3194_ _3431_/CLK _3194_/D vssd1 vssd1 vccd1 vccd1 _3194_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2145_ _3350_/Q _2146_/B vssd1 vssd1 vccd1 vccd1 _2152_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_88_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2076_ _2092_/A _2059_/Y _2060_/Y _2058_/C vssd1 vssd1 vccd1 vccd1 _2076_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1642__A1 _2576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2978_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2978_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1929_ _1929_/A _1929_/B vssd1 vssd1 vccd1 vccd1 _1930_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_71_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold730 _3193_/Q vssd1 vssd1 vccd1 vccd1 hold730/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold752 _3174_/Q vssd1 vssd1 vccd1 vccd1 hold752/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 _2617_/X vssd1 vssd1 vccd1 vccd1 _3165_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 _2909_/X vssd1 vssd1 vccd1 vccd1 _3437_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 _3512_/Q vssd1 vssd1 vccd1 vccd1 _2349_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold796 _3505_/Q vssd1 vssd1 vccd1 vccd1 hold796/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 _2022_/X vssd1 vssd1 vccd1 vccd1 _3504_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1633__S hold12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2658__A0 _2801_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1633__A1 hold59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2649__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2901_ _2901_/A _2901_/B vssd1 vssd1 vccd1 vccd1 _2910_/S sky130_fd_sc_hd__nand2_4
X_2832_ _2098_/S hold560/X _2839_/S vssd1 vssd1 vccd1 vccd1 _2832_/X sky130_fd_sc_hd__mux2_1
X_2763_ _2803_/A1 hold341/X _2769_/S vssd1 vssd1 vccd1 vccd1 _2763_/X sky130_fd_sc_hd__mux2_1
X_1714_ _3536_/Q _3453_/Q vssd1 vssd1 vccd1 vccd1 _1714_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_5_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2403__A hold70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2694_ hold394/X _2806_/A1 _2697_/S vssd1 vssd1 vccd1 vccd1 _2694_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1645_ _2289_/A hold52/X vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__nor2_1
X_1576_ _3605_/Q vssd1 vssd1 vccd1 vccd1 _1576_/Y sky130_fd_sc_hd__inv_2
X_3315_ _3324_/CLK hold39/X vssd1 vssd1 vccd1 vccd1 _3315_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ _3318_/CLK _3246_/D vssd1 vssd1 vccd1 vccd1 _3246_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3177_ _3619_/CLK _3177_/D vssd1 vssd1 vccd1 vccd1 _3177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2128_ _2379_/C _2377_/C vssd1 vssd1 vccd1 vccd1 _2133_/B sky130_fd_sc_hd__nand2_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2059_ _3546_/Q _2084_/B vssd1 vssd1 vccd1 vccd1 _2059_/Y sky130_fd_sc_hd__nand2_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold560 _3363_/Q vssd1 vssd1 vccd1 vccd1 hold560/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold571 _2814_/X vssd1 vssd1 vccd1 vccd1 _3337_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2879__A0 _2355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold582 _3433_/Q vssd1 vssd1 vccd1 vccd1 hold582/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 _2908_/X vssd1 vssd1 vccd1 vccd1 _3436_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1765__C _1769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3100_ _3101_/A vssd1 vssd1 vccd1 vccd1 _3100_/Y sky130_fd_sc_hd__inv_2
X_3031_ _3032_/A vssd1 vssd1 vccd1 vccd1 _3031_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_3_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3509_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2815_ hold536/X _2104_/B _2819_/S vssd1 vssd1 vccd1 vccd1 _2815_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2746_ _2806_/A1 hold273/X _2749_/S vssd1 vssd1 vccd1 vccd1 _2746_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2677_ _3488_/Q _2677_/B hold36/X vssd1 vssd1 vccd1 vccd1 _2760_/A sky130_fd_sc_hd__or3b_2
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1628_ _2289_/A hold11/X vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__nor2_1
X_1559_ _3630_/Q vssd1 vssd1 vccd1 vccd1 _1559_/Y sky130_fd_sc_hd__inv_2
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3229_ _3326_/CLK _3229_/D vssd1 vssd1 vccd1 vccd1 _3229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2742__S _2749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2978__A _3124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold390 _3600_/Q vssd1 vssd1 vccd1 vccd1 hold390/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2652__S _2654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3580_ _3590_/CLK _3580_/D _3071_/Y vssd1 vssd1 vccd1 vccd1 _3580_/Q sky130_fd_sc_hd__dfrtp_1
X_2600_ _2355_/B hold700/X _2601_/S vssd1 vssd1 vccd1 vccd1 _2600_/X sky130_fd_sc_hd__mux2_1
X_2531_ _3378_/Q _3360_/Q _3369_/Q _3197_/Q _1918_/B _1912_/B vssd1 vssd1 vccd1 vccd1
+ _2531_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2307__A2 _2064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2462_ _3442_/Q hold21/A _2461_/X _2574_/A vssd1 vssd1 vccd1 vccd1 _2462_/X sky130_fd_sc_hd__o211a_1
X_2393_ _3593_/Q _3384_/Q _3344_/Q _3595_/Q _2390_/X vssd1 vssd1 vccd1 vccd1 _2395_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2827__S _2829_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3014_ _3110_/A vssd1 vssd1 vccd1 vccd1 _3014_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1967__A _2144_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2729_ _2708_/A _2729_/B vssd1 vssd1 vccd1 vccd1 _2760_/B sky130_fd_sc_hd__nand2b_2
Xfanout122 input2/X vssd1 vssd1 vccd1 vccd1 _3097_/A sky130_fd_sc_hd__buf_8
Xfanout100 hold994/X vssd1 vssd1 vccd1 vccd1 _1811_/S sky130_fd_sc_hd__clkbuf_4
Xfanout111 hold126/X vssd1 vssd1 vccd1 vccd1 _2399_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1641__S hold12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2220__B _2221_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2647__S _2654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1962_ _3297_/Q hold42/X hold349/X hold343/X _2049_/S0 _2195_/A1 vssd1 vssd1 vccd1
+ vccd1 _1962_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_83_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1893_ _2613_/B _1893_/B vssd1 vssd1 vccd1 vccd1 _1893_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3632_ _3632_/CLK hold16/X _3123_/Y vssd1 vssd1 vccd1 vccd1 _3632_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3563_ _3567_/CLK _3563_/D _3057_/Y vssd1 vssd1 vccd1 vccd1 _3563_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2514_ _2574_/A _2505_/X _2506_/X _2513_/X vssd1 vssd1 vccd1 vccd1 _2514_/X sky130_fd_sc_hd__o22a_2
X_3494_ _3635_/CLK _3494_/D _2988_/Y vssd1 vssd1 vccd1 vccd1 _3494_/Q sky130_fd_sc_hd__dfrtp_1
X_2445_ _3441_/Q hold21/A _2444_/X _2574_/A vssd1 vssd1 vccd1 vccd1 _2445_/X sky130_fd_sc_hd__o211a_1
X_2376_ _1793_/B _1826_/Y _2370_/A _1769_/B _1808_/D vssd1 vssd1 vccd1 vccd1 _2376_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_78_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1636__S hold12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _2230_/A _2230_/B vssd1 vssd1 vccd1 vccd1 _2234_/A sky130_fd_sc_hd__nand2_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2694__A1 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2161_ _1945_/A _2161_/B _2161_/C _2161_/D vssd1 vssd1 vccd1 vccd1 _2162_/C sky130_fd_sc_hd__and4b_1
XFILLER_0_88_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2092_ _2092_/A _3539_/Q vssd1 vssd1 vccd1 vccd1 _2092_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2541__S1 _1912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2994_ _3057_/A vssd1 vssd1 vccd1 vccd1 _2994_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2406__A _2406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1945_ _1945_/A _2161_/B vssd1 vssd1 vccd1 vccd1 _1945_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1876_ _1837_/A _1844_/Y _1875_/X _1843_/A _1836_/A vssd1 vssd1 vccd1 vccd1 _1876_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold912 _3500_/Q vssd1 vssd1 vccd1 vccd1 _1588_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3615_ _3627_/CLK hold76/X _3106_/Y vssd1 vssd1 vccd1 vccd1 _3615_/Q sky130_fd_sc_hd__dfrtp_1
Xhold901 _3149_/Q vssd1 vssd1 vccd1 vccd1 _1808_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 _3533_/Q vssd1 vssd1 vccd1 vccd1 _1865_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold945 _1752_/X vssd1 vssd1 vccd1 vccd1 _3564_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3546_ _3555_/CLK _3546_/D _3040_/Y vssd1 vssd1 vccd1 vccd1 _3546_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout104_A hold70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold934 _2142_/Y vssd1 vssd1 vccd1 vccd1 _2143_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 _2233_/X vssd1 vssd1 vccd1 vccd1 _2234_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 _1750_/X vssd1 vssd1 vccd1 vccd1 _3565_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 _3562_/Q vssd1 vssd1 vccd1 vccd1 _1753_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 _1823_/Y vssd1 vssd1 vccd1 vccd1 _1824_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3477_ _3533_/CLK _3477_/D _2971_/Y vssd1 vssd1 vccd1 vccd1 _3477_/Q sky130_fd_sc_hd__dfrtp_1
X_2428_ _3181_/Q _3334_/Q _3163_/Q _3139_/Q _1944_/B _1943_/A vssd1 vssd1 vccd1 vccd1
+ _2428_/X sky130_fd_sc_hd__mux4_1
X_2359_ _3616_/Q _2360_/B vssd1 vssd1 vccd1 vccd1 _2359_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2532__S1 _2532_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2676__A1 _2406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1730_ _3531_/Q _1730_/B vssd1 vssd1 vccd1 vccd1 _1730_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_80_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1661_ hold98/A _1661_/B _2416_/A vssd1 vssd1 vccd1 vccd1 _1661_/X sky130_fd_sc_hd__and3_1
Xhold208 _3233_/Q vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 _2717_/X vssd1 vssd1 vccd1 vccd1 _3251_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3057__A _3057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3400_ _3521_/CLK _3400_/D vssd1 vssd1 vccd1 vccd1 _3400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2364__B1 _2109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3331_ _3509_/CLK _3331_/D vssd1 vssd1 vccd1 vccd1 _3331_/Q sky130_fd_sc_hd__dfxtp_1
X_1592_ _1957_/A vssd1 vssd1 vccd1 vccd1 _2184_/A sky130_fd_sc_hd__inv_2
XFILLER_0_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3321_/CLK _3262_/D vssd1 vssd1 vccd1 vccd1 _3262_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ _2213_/A _2213_/B vssd1 vssd1 vccd1 vccd1 _2213_/X sky130_fd_sc_hd__or2_1
X_3193_ _3424_/CLK _3193_/D vssd1 vssd1 vccd1 vccd1 _3193_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2144_ _2144_/A _2379_/A _2144_/C _2144_/D vssd1 vssd1 vccd1 vccd1 _2146_/B sky130_fd_sc_hd__or4_1
X_2075_ _2356_/B _2075_/B vssd1 vssd1 vccd1 vccd1 _2099_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2977_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2977_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1928_ _2349_/B _1929_/B _1927_/Y vssd1 vssd1 vccd1 vccd1 _1931_/A sky130_fd_sc_hd__a21bo_1
X_1859_ _1859_/A _1859_/B vssd1 vssd1 vccd1 vccd1 _1859_/X sky130_fd_sc_hd__or2_1
Xhold720 _3391_/Q vssd1 vssd1 vccd1 vccd1 hold720/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold753 _2627_/X vssd1 vssd1 vccd1 vccd1 _3174_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 _3366_/Q vssd1 vssd1 vccd1 vccd1 hold764/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 _2649_/X vssd1 vssd1 vccd1 vccd1 _3193_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 _3390_/Q vssd1 vssd1 vccd1 vccd1 hold742/X sky130_fd_sc_hd__dlygate4sd3_1
X_3529_ _3532_/CLK _3529_/D _3023_/Y vssd1 vssd1 vccd1 vccd1 _3529_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2450__S0 _2532_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold786 hold786/A vssd1 vssd1 vccd1 vccd1 _1708_/B sky130_fd_sc_hd__buf_1
Xhold775 _1940_/X vssd1 vssd1 vccd1 vccd1 _3512_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 _2012_/X vssd1 vssd1 vccd1 vccd1 _3505_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2745__S _2749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_27_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3559_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_35_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2594__A0 _2098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
X_2900_ hold490/X _2058_/X _2900_/S vssd1 vssd1 vccd1 vccd1 _2900_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2821__A1 _2358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2831_ _2358_/B hold768/X _2839_/S vssd1 vssd1 vccd1 vccd1 _2831_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2762_ _2802_/A1 hold142/X _2769_/S vssd1 vssd1 vccd1 vccd1 _2762_/X sky130_fd_sc_hd__mux2_1
X_1713_ _1724_/B _1883_/A vssd1 vssd1 vccd1 vccd1 _1713_/Y sky130_fd_sc_hd__nand2b_1
X_2693_ hold397/X _2805_/A1 _2697_/S vssd1 vssd1 vccd1 vccd1 _2693_/X sky130_fd_sc_hd__mux2_1
X_1644_ hold51/X _1644_/B vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__or2_2
X_1575_ _3606_/Q vssd1 vssd1 vccd1 vccd1 _1575_/Y sky130_fd_sc_hd__inv_2
X_3314_ _3324_/CLK _3314_/D vssd1 vssd1 vccd1 vccd1 _3314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _3319_/CLK _3245_/D vssd1 vssd1 vccd1 vccd1 _3245_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3176_ _3424_/CLK _3176_/D vssd1 vssd1 vccd1 vccd1 _3176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2127_ _2127_/A _2127_/B _2127_/C _2127_/D vssd1 vssd1 vccd1 vccd1 _2377_/C sky130_fd_sc_hd__and4_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2058_ _2063_/A _2096_/B _2058_/C _2058_/D vssd1 vssd1 vccd1 vccd1 _2058_/X sky130_fd_sc_hd__and4bb_2
XFILLER_0_88_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2499__S0 _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2812__A1 _2098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold550 _3413_/Q vssd1 vssd1 vccd1 vccd1 hold550/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 _2832_/X vssd1 vssd1 vccd1 vccd1 _3363_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 _3186_/Q vssd1 vssd1 vccd1 vccd1 hold572/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 _2905_/X vssd1 vssd1 vccd1 vccd1 _3433_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 _3139_/Q vssd1 vssd1 vccd1 vccd1 hold594/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout84_A _2532_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2803__A1 _2803_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output65_A _2540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3030_ _3032_/A vssd1 vssd1 vccd1 vccd1 _3030_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2814_ hold570/X _2105_/A _2819_/S vssd1 vssd1 vccd1 vccd1 _2814_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2745_ _2805_/A1 hold297/X _2749_/S vssd1 vssd1 vccd1 vccd1 _2745_/X sky130_fd_sc_hd__mux2_1
X_2676_ hold433/X _2406_/A _2676_/S vssd1 vssd1 vccd1 vccd1 _2676_/X sky130_fd_sc_hd__mux2_1
X_1627_ hold9/X _1644_/B vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__or2_1
XFILLER_0_1_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1558_ hold27/X vssd1 vssd1 vccd1 vccd1 _1558_/Y sky130_fd_sc_hd__inv_2
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3228_ _3320_/CLK _3228_/D vssd1 vssd1 vccd1 vccd1 _3228_/Q sky130_fd_sc_hd__dfxtp_1
X_3159_ _3619_/CLK _3159_/D vssd1 vssd1 vccd1 vccd1 _3159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1639__S hold12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold380 _3322_/Q vssd1 vssd1 vccd1 vccd1 hold380/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2721__A0 _2802_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold391 _3613_/Q vssd1 vssd1 vccd1 vccd1 _1569_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2994__A _3057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_42_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3516_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2788__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2530_ _2529_/X _2528_/X _2546_/S vssd1 vssd1 vccd1 vccd1 _2530_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2461_ _3636_/Q _2510_/A _2458_/X _2460_/X _2510_/B vssd1 vssd1 vccd1 vccd1 _2461_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2712__A0 _2803_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2392_ hold68/A _3381_/Q _3346_/Q hold85/A vssd1 vssd1 vccd1 vccd1 _2392_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_64_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3013_ _3110_/A vssd1 vssd1 vccd1 vccd1 _3013_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2843__S _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2728_ _2406_/A hold403/X _2728_/S vssd1 vssd1 vccd1 vccd1 _2728_/X sky130_fd_sc_hd__mux2_1
X_2659_ _2802_/A1 hold171/X _2666_/S vssd1 vssd1 vccd1 vccd1 _2659_/X sky130_fd_sc_hd__mux2_1
Xfanout112 hold123/X vssd1 vssd1 vccd1 vccd1 _2801_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__2703__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout101 hold30/X vssd1 vssd1 vccd1 vccd1 _2406_/A sky130_fd_sc_hd__clkbuf_8
Xfanout123 _3124_/A vssd1 vssd1 vccd1 vccd1 _3122_/A sky130_fd_sc_hd__buf_8
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1961_ _1959_/X _1960_/X _2036_/S vssd1 vssd1 vccd1 vccd1 _1961_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1892_ _1892_/A _1896_/A vssd1 vssd1 vccd1 vccd1 _1893_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3631_ _3633_/CLK hold81/X _3122_/Y vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__dfstp_1
XFILLER_0_36_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3562_ _3567_/CLK _3562_/D _3056_/Y vssd1 vssd1 vccd1 vccd1 _3562_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2513_ _3625_/Q hold11/A _2559_/B _2512_/X vssd1 vssd1 vccd1 vccd1 _2513_/X sky130_fd_sc_hd__o211a_1
X_3493_ _3576_/CLK _3493_/D _2987_/Y vssd1 vssd1 vccd1 vccd1 _3493_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2444_ _3635_/Q _2510_/A _2441_/X _2443_/X _2510_/B vssd1 vssd1 vccd1 vccd1 _2444_/X
+ sky130_fd_sc_hd__a221o_1
X_2375_ _2375_/A _2375_/B vssd1 vssd1 vccd1 vccd1 _3347_/D sky130_fd_sc_hd__nand2_1
XANTENNA__1672__A0 _2576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2748__S _2749_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ _3521_/Q _2160_/B vssd1 vssd1 vccd1 vccd1 _2161_/D sky130_fd_sc_hd__xnor2_1
X_2091_ _2080_/Y _2083_/Y _2091_/S vssd1 vssd1 vccd1 vccd1 _2091_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2993_ _3129_/A vssd1 vssd1 vccd1 vccd1 _2993_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_61_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1944_ _3519_/Q _1944_/B vssd1 vssd1 vccd1 vccd1 _2161_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1875_ _3527_/Q _1877_/B _1843_/A vssd1 vssd1 vccd1 vccd1 _1875_/X sky130_fd_sc_hd__a21o_1
X_3614_ _3614_/CLK _3614_/D _3105_/Y vssd1 vssd1 vccd1 vccd1 _3614_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2906__A0 _2104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold902 _2374_/X vssd1 vssd1 vccd1 vccd1 _3149_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 _2118_/Y vssd1 vssd1 vccd1 vccd1 _3500_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 _3535_/Q vssd1 vssd1 vccd1 vccd1 _1851_/A sky130_fd_sc_hd__buf_1
Xhold924 _1866_/X vssd1 vssd1 vccd1 vccd1 _3533_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3545_ _3571_/CLK _3545_/D _3039_/Y vssd1 vssd1 vccd1 vccd1 _3545_/Q sky130_fd_sc_hd__dfrtp_1
Xhold935 _2143_/Y vssd1 vssd1 vccd1 vccd1 _3496_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3476_ _3533_/CLK _3476_/D _2970_/Y vssd1 vssd1 vccd1 vccd1 _3476_/Q sky130_fd_sc_hd__dfrtp_1
Xhold979 _3563_/Q vssd1 vssd1 vccd1 vccd1 hold979/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 _1756_/X vssd1 vssd1 vccd1 vccd1 _3562_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 _3557_/Q vssd1 vssd1 vccd1 vccd1 hold957/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2382__A1 _2000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2427_ _3403_/Q _3394_/Q _3385_/Q _3430_/Q _1944_/B _1943_/A vssd1 vssd1 vccd1 vccd1
+ _2427_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_86_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2134__A1 _2000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2358_ _2358_/A _2358_/B vssd1 vssd1 vccd1 vccd1 _2367_/D sky130_fd_sc_hd__xnor2_1
X_2289_ _2289_/A hold21/X vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__nor2_2
XFILLER_0_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1948__A1 _3518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2048__S1 _2219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1890__B _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1660_ _2165_/B _2421_/A vssd1 vssd1 vccd1 vccd1 _2435_/A sky130_fd_sc_hd__and2_2
X_1591_ _2228_/C vssd1 vssd1 vccd1 vccd1 _1591_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold209 _2696_/X vssd1 vssd1 vccd1 vccd1 _3233_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3330_ _3330_/CLK _3330_/D vssd1 vssd1 vccd1 vccd1 _3330_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _3333_/CLK _3261_/D vssd1 vssd1 vccd1 vccd1 _3261_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ _2209_/X _2210_/Y _2211_/Y _2211_/B _2208_/A vssd1 vssd1 vccd1 vccd1 _2212_/X
+ sky130_fd_sc_hd__a32o_1
X_3192_ _3413_/CLK _3192_/D vssd1 vssd1 vccd1 vccd1 _3192_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2143_ _2143_/A _2143_/B vssd1 vssd1 vccd1 vccd1 _2143_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__1970__S0 _3483_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2074_ _2061_/X _2357_/B _2355_/B _2071_/X vssd1 vssd1 vccd1 vccd1 _2075_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_88_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2976_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2976_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1927_ _1941_/S _1939_/B vssd1 vssd1 vccd1 vccd1 _1927_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1858_ _1858_/A _1858_/B vssd1 vssd1 vccd1 vccd1 _3537_/D sky130_fd_sc_hd__and2_1
Xhold710 _3141_/Q vssd1 vssd1 vccd1 vccd1 hold710/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 _2858_/X vssd1 vssd1 vccd1 vccd1 _3391_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 _3370_/Q vssd1 vssd1 vccd1 vccd1 hold732/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 _3388_/Q vssd1 vssd1 vccd1 vccd1 hold754/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold743 _2857_/X vssd1 vssd1 vccd1 vccd1 _3390_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1789_ _2319_/A _2308_/B vssd1 vssd1 vccd1 vccd1 _2126_/B sky130_fd_sc_hd__nor2_1
X_3528_ _3532_/CLK _3528_/D _3022_/Y vssd1 vssd1 vccd1 vccd1 _3528_/Q sky130_fd_sc_hd__dfrtp_1
Xhold765 _2835_/X vssd1 vssd1 vccd1 vccd1 _3366_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2450__S1 _1912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold776 _3376_/Q vssd1 vssd1 vccd1 vccd1 hold776/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 _1708_/X vssd1 vssd1 vccd1 vccd1 _3568_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3459_ _3594_/CLK _3459_/D _2953_/Y vssd1 vssd1 vccd1 vccd1 _3459_/Q sky130_fd_sc_hd__dfrtp_1
Xhold798 _3465_/Q vssd1 vssd1 vccd1 vccd1 _2249_/A sky130_fd_sc_hd__buf_1
XANTENNA__2107__B2 _2064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1618__A0 _1767_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2291__A0 _3454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2761__S _2769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2001__S _2055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__buf_2
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2830_ _2881_/B _2830_/B vssd1 vssd1 vccd1 vccd1 _2839_/S sky130_fd_sc_hd__nand2_4
XFILLER_0_42_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2761_ _2801_/A1 hold288/X _2769_/S vssd1 vssd1 vccd1 vccd1 _2761_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1712_ _3454_/Q _1853_/A vssd1 vssd1 vccd1 vccd1 _1712_/X sky130_fd_sc_hd__and2b_1
XANTENNA__2585__A1 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2692_ hold206/X _2804_/A1 _2697_/S vssd1 vssd1 vccd1 vccd1 _2692_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1643_ hold93/A _1644_/B vssd1 vssd1 vccd1 vccd1 _1643_/Y sky130_fd_sc_hd__nor2_2
X_1574_ _1574_/A vssd1 vssd1 vccd1 vccd1 _1574_/Y sky130_fd_sc_hd__inv_2
X_3313_ _3322_/CLK _3313_/D vssd1 vssd1 vccd1 vccd1 _3313_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _3321_/CLK _3244_/D vssd1 vssd1 vccd1 vccd1 _3244_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2846__S _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3175_ _3424_/CLK _3175_/D vssd1 vssd1 vccd1 vccd1 _3175_/Q sky130_fd_sc_hd__dfxtp_1
X_2126_ _2126_/A _2126_/B vssd1 vssd1 vccd1 vccd1 _2127_/D sky130_fd_sc_hd__nand2_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2057_ _2121_/A _3547_/Q _2084_/B vssd1 vssd1 vccd1 vccd1 _2096_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_88_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2499__S1 _1943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2581__S _2589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2959_ _3069_/A vssd1 vssd1 vccd1 vccd1 _2959_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold551 _2883_/X vssd1 vssd1 vccd1 vccd1 _3413_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold540 _3192_/Q vssd1 vssd1 vccd1 vccd1 hold540/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 _3142_/Q vssd1 vssd1 vccd1 vccd1 hold562/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold595 _2593_/X vssd1 vssd1 vccd1 vccd1 _3139_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold584 _3342_/Q vssd1 vssd1 vccd1 vccd1 hold584/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 _2640_/X vssd1 vssd1 vccd1 vccd1 _3186_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput60 _3655_/A vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_12
X_2813_ hold588/X _2109_/B _2819_/S vssd1 vssd1 vccd1 vccd1 _2813_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2744_ _2804_/A1 hold159/X _2749_/S vssd1 vssd1 vccd1 vccd1 _2744_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2675_ hold319/X _2808_/A1 _2676_/S vssd1 vssd1 vccd1 vccd1 _2675_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1626_ hold35/X _1626_/B vssd1 vssd1 vccd1 vccd1 _1644_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1557_ _1557_/A vssd1 vssd1 vccd1 vccd1 _1836_/A sky130_fd_sc_hd__clkinv_4
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3227_ _3408_/CLK _3227_/D vssd1 vssd1 vccd1 vccd1 _3227_/Q sky130_fd_sc_hd__dfxtp_1
X_3158_ _3431_/CLK _3158_/D vssd1 vssd1 vccd1 vccd1 _3158_/Q sky130_fd_sc_hd__dfxtp_1
X_2109_ _2360_/B _2109_/B vssd1 vssd1 vccd1 vccd1 _2110_/B sky130_fd_sc_hd__xor2_1
X_3089_ _3090_/A vssd1 vssd1 vccd1 vccd1 _3089_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_64_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2797__A1 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold370 _3277_/Q vssd1 vssd1 vccd1 vccd1 hold370/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 _2797_/X vssd1 vssd1 vccd1 vccd1 _3322_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 _3240_/Q vssd1 vssd1 vccd1 vccd1 hold392/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2486__S _3518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_11_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3321_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2460_ _3622_/Q hold11/A hold52/A _3613_/Q _2459_/X vssd1 vssd1 vccd1 vccd1 _2460_/X
+ sky130_fd_sc_hd__o221a_1
X_2391_ _3592_/Q _3590_/Q _3380_/Q _3598_/Q vssd1 vssd1 vccd1 vccd1 _2395_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3012_ _3110_/A vssd1 vssd1 vccd1 vccd1 _3012_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2779__A1 hold30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout127_A _3057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2727_ _2808_/A1 hold196/X _2728_/S vssd1 vssd1 vccd1 vccd1 _2727_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2658_ _2801_/A1 hold290/X _2666_/S vssd1 vssd1 vccd1 vccd1 _2658_/X sky130_fd_sc_hd__mux2_1
X_1609_ input6/X input7/X hold33/X input9/X vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__or4_1
X_2589_ hold409/X _2406_/A _2589_/S vssd1 vssd1 vccd1 vccd1 _2589_/X sky130_fd_sc_hd__mux2_1
Xfanout102 hold45/X vssd1 vssd1 vccd1 vccd1 _2808_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout113 hold123/X vssd1 vssd1 vccd1 vccd1 _2576_/A sky130_fd_sc_hd__clkbuf_4
Xfanout124 input2/X vssd1 vssd1 vccd1 vccd1 _3124_/A sky130_fd_sc_hd__buf_8
XFILLER_0_77_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1681__A1 hold87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1960_ hold425/X hold433/X hold399/X hold413/X _2045_/S0 _2045_/S1 vssd1 vssd1 vccd1
+ vccd1 _1960_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2630__A0 _2360_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1891_ _1891_/A _1902_/A _3519_/Q vssd1 vssd1 vccd1 vccd1 _1896_/A sky130_fd_sc_hd__and3_1
XFILLER_0_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3630_ _3633_/CLK hold13/X _3121_/Y vssd1 vssd1 vccd1 vccd1 _3630_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_70_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3561_ _3567_/CLK _3561_/D _3055_/Y vssd1 vssd1 vccd1 vccd1 _3561_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2512_ _3616_/Q _1643_/Y _2572_/C _2511_/X vssd1 vssd1 vccd1 vccd1 _2512_/X sky130_fd_sc_hd__a22o_1
X_3492_ _3576_/CLK _3492_/D _2986_/Y vssd1 vssd1 vccd1 vccd1 _3492_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2443_ _2070_/A hold11/A hold52/A _3612_/Q _2442_/X vssd1 vssd1 vccd1 vccd1 _2443_/X
+ sky130_fd_sc_hd__o221a_1
X_2374_ _1808_/B _2373_/X _2387_/C vssd1 vssd1 vccd1 vccd1 _2374_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2544__S0 _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2621__A0 _2357_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2764__S _2769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2860__A0 _2356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1663__A1 _2400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2612__A0 _2356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2679__A0 _2801_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output40_A _3577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2090_ _2090_/A _2090_/B vssd1 vssd1 vccd1 vccd1 _2095_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1654__A1 _2576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2992_ _3049_/A vssd1 vssd1 vccd1 vccd1 _2992_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_83_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1943_ _1943_/A _1943_/B vssd1 vssd1 vccd1 vccd1 _1945_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1874_ _1873_/Y _1871_/B _1845_/A _1836_/A vssd1 vssd1 vccd1 vccd1 _3529_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_71_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3613_ _3614_/CLK _3613_/D _3104_/Y vssd1 vssd1 vccd1 vccd1 _3613_/Q sky130_fd_sc_hd__dfrtp_1
Xhold903 _3348_/Q vssd1 vssd1 vccd1 vccd1 _2379_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 _3530_/Q vssd1 vssd1 vccd1 vccd1 _1871_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold936 _3524_/Q vssd1 vssd1 vccd1 vccd1 _1883_/A sky130_fd_sc_hd__clkbuf_2
Xhold914 _3486_/Q vssd1 vssd1 vccd1 vccd1 hold914/X sky130_fd_sc_hd__dlygate4sd3_1
X_3544_ _3573_/CLK _3544_/D _3038_/Y vssd1 vssd1 vccd1 vccd1 _3544_/Q sky130_fd_sc_hd__dfrtp_1
Xhold947 _1862_/X vssd1 vssd1 vccd1 vccd1 _3535_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3475_ _3532_/CLK _3475_/D _2969_/Y vssd1 vssd1 vccd1 vccd1 _3475_/Q sky130_fd_sc_hd__dfrtp_1
Xhold969 _3559_/Q vssd1 vssd1 vccd1 vccd1 hold969/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 _1766_/X vssd1 vssd1 vccd1 vccd1 _3557_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2849__S _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2426_ _3440_/Q hold21/A _2425_/X _2574_/A vssd1 vssd1 vccd1 vccd1 _2426_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_86_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2357_ hold90/X _2357_/B vssd1 vssd1 vccd1 vccd1 _2363_/D sky130_fd_sc_hd__xnor2_1
X_2288_ hold35/X hold20/X vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__nand2_2
XANTENNA__2584__S _2589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2833__A0 _2109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1636__A1 hold87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1590_ _2221_/B vssd1 vssd1 vccd1 vccd1 _2193_/A sky130_fd_sc_hd__inv_2
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2364__A2 _2098_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _3332_/CLK _3260_/D vssd1 vssd1 vccd1 vccd1 _3260_/Q sky130_fd_sc_hd__dfxtp_1
X_2211_ _2211_/A _2211_/B vssd1 vssd1 vccd1 vccd1 _2211_/Y sky130_fd_sc_hd__nor2_1
X_3191_ _3413_/CLK _3191_/D vssd1 vssd1 vccd1 vccd1 _3191_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2142_ _2130_/A _2139_/B _2139_/A vssd1 vssd1 vccd1 vccd1 _2142_/Y sky130_fd_sc_hd__a21oi_1
X_2073_ _2061_/X _2106_/B vssd1 vssd1 vccd1 vccd1 _2073_/X sky130_fd_sc_hd__and2b_1
XANTENNA__1970__S1 _2045_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2975_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2975_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1926_ _2349_/B _1932_/B vssd1 vssd1 vccd1 vccd1 _1939_/B sky130_fd_sc_hd__xor2_1
X_1857_ _1859_/A _1837_/A _1859_/B _1853_/A vssd1 vssd1 vccd1 vccd1 _1858_/B sky130_fd_sc_hd__a31o_1
Xhold700 _3146_/Q vssd1 vssd1 vccd1 vccd1 hold700/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold711 _2595_/X vssd1 vssd1 vccd1 vccd1 _3141_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3527_ _3532_/CLK _3527_/D _3021_/Y vssd1 vssd1 vccd1 vccd1 _3527_/Q sky130_fd_sc_hd__dfrtp_1
Xhold744 _3412_/Q vssd1 vssd1 vccd1 vccd1 hold744/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 _2839_/X vssd1 vssd1 vccd1 vccd1 _3370_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 _2855_/X vssd1 vssd1 vccd1 vccd1 _3388_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 _3154_/Q vssd1 vssd1 vccd1 vccd1 hold722/X sky130_fd_sc_hd__dlygate4sd3_1
X_1788_ _2091_/S _2064_/A _1564_/Y vssd1 vssd1 vccd1 vccd1 _2308_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_12_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold766 _3158_/Q vssd1 vssd1 vccd1 vccd1 hold766/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 _2846_/X vssd1 vssd1 vccd1 vccd1 _3376_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 _3508_/Q vssd1 vssd1 vccd1 vccd1 hold788/X sky130_fd_sc_hd__dlygate4sd3_1
X_3458_ _3594_/CLK _3458_/D _2952_/Y vssd1 vssd1 vccd1 vccd1 _3458_/Q sky130_fd_sc_hd__dfrtp_1
Xhold799 _2255_/X vssd1 vssd1 vccd1 vccd1 _3466_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3389_ _3434_/CLK _3389_/D vssd1 vssd1 vccd1 vccd1 _3389_/Q sky130_fd_sc_hd__dfxtp_1
X_2409_ _2438_/B vssd1 vssd1 vccd1 vccd1 _2409_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1618__A1 hold75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2043__A1 _2144_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3575_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2760_ _2760_/A _2760_/B vssd1 vssd1 vccd1 vccd1 _2769_/S sky130_fd_sc_hd__or2_4
X_1711_ _3455_/Q _1855_/A vssd1 vssd1 vccd1 vccd1 _1711_/Y sky130_fd_sc_hd__nand2b_1
X_2691_ hold324/X _2803_/A1 _2697_/S vssd1 vssd1 vccd1 vccd1 _2691_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1642_ _2121_/A _2576_/A hold12/X vssd1 vssd1 vccd1 vccd1 _3620_/D sky130_fd_sc_hd__mux2_1
XANTENNA__2337__A2 _2363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1573_ _1573_/A vssd1 vssd1 vccd1 vccd1 _2349_/A sky130_fd_sc_hd__inv_2
X_3312_ _3321_/CLK _3312_/D vssd1 vssd1 vccd1 vccd1 _3312_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _3408_/CLK _3243_/D vssd1 vssd1 vccd1 vccd1 _3243_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ _3579_/CLK _3174_/D vssd1 vssd1 vccd1 vccd1 _3174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2125_ _2126_/A _2126_/B vssd1 vssd1 vccd1 vccd1 _2127_/C sky130_fd_sc_hd__or2_1
XFILLER_0_88_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2056_ _2063_/A _2070_/A _2058_/D vssd1 vssd1 vccd1 vccd1 _2084_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__2862__S _2870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2958_ _3069_/A vssd1 vssd1 vccd1 vccd1 _2958_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1909_ _1922_/A _2871_/C vssd1 vssd1 vccd1 vccd1 _1909_/Y sky130_fd_sc_hd__nand2_1
X_2889_ _2073_/X hold566/X _2890_/S vssd1 vssd1 vccd1 vccd1 _2889_/X sky130_fd_sc_hd__mux2_1
Xhold530 _3422_/Q vssd1 vssd1 vccd1 vccd1 hold530/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold541 _2648_/X vssd1 vssd1 vccd1 vccd1 _3192_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 _3374_/Q vssd1 vssd1 vccd1 vccd1 hold552/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 _2596_/X vssd1 vssd1 vccd1 vccd1 _3142_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 _3414_/Q vssd1 vssd1 vccd1 vccd1 hold596/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 _2819_/X vssd1 vssd1 vccd1 vccd1 _3342_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 _3144_/Q vssd1 vssd1 vccd1 vccd1 hold574/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2772__S _2779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput61 _2487_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_12
Xoutput50 _3648_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_12
XANTENNA__2012__S _2055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2812_ hold548/X _2098_/S _2819_/S vssd1 vssd1 vccd1 vccd1 _2812_/X sky130_fd_sc_hd__mux2_1
X_2743_ _2803_/A1 hold347/X _2749_/S vssd1 vssd1 vccd1 vccd1 _2743_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2674_ hold429/X _2807_/A1 _2676_/S vssd1 vssd1 vccd1 vccd1 _2674_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1625_ _1625_/A vssd1 vssd1 vccd1 vccd1 _1626_/B sky130_fd_sc_hd__inv_2
XFILLER_0_1_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1556_ _1950_/A vssd1 vssd1 vccd1 vccd1 _2381_/A sky130_fd_sc_hd__inv_2
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3226_ _3320_/CLK _3226_/D vssd1 vssd1 vccd1 vccd1 _3226_/Q sky130_fd_sc_hd__dfxtp_1
X_3157_ _3424_/CLK _3157_/D vssd1 vssd1 vccd1 vccd1 _3157_/Q sky130_fd_sc_hd__dfxtp_1
X_2108_ _2090_/A _2071_/X _2107_/X vssd1 vssd1 vccd1 vccd1 _2108_/Y sky130_fd_sc_hd__a21oi_2
X_3088_ _3090_/A vssd1 vssd1 vccd1 vccd1 _3088_/Y sky130_fd_sc_hd__inv_2
X_2039_ _2038_/X _2037_/X _2222_/A vssd1 vssd1 vccd1 vccd1 _2040_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_9_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold371 _2747_/X vssd1 vssd1 vccd1 vccd1 _3277_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold360 _2716_/X vssd1 vssd1 vccd1 vccd1 _3250_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2767__S _2769_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold393 _2704_/X vssd1 vssd1 vccd1 vccd1 _3240_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _3327_/Q vssd1 vssd1 vccd1 vccd1 hold382/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2007__S _2036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_51_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3438_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2390_ _3600_/Q _3382_/Q _3343_/Q hold82/A vssd1 vssd1 vccd1 vccd1 _2390_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3011_ _3110_/A vssd1 vssd1 vccd1 vccd1 _3011_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_64_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1610__A _1657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2144__C _2144_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2726_ _2807_/A1 hold401/X _2728_/S vssd1 vssd1 vccd1 vccd1 _2726_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2657_ hold37/X _2800_/B vssd1 vssd1 vccd1 vccd1 _2666_/S sky130_fd_sc_hd__or2_4
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1608_ _1608_/A _2577_/B vssd1 vssd1 vccd1 vccd1 _2289_/A sky130_fd_sc_hd__nand2_2
Xfanout103 hold87/X vssd1 vssd1 vccd1 vccd1 _2807_/A1 sky130_fd_sc_hd__buf_4
X_2588_ hold222/X _2808_/A1 _2589_/S vssd1 vssd1 vccd1 vccd1 _2588_/X sky130_fd_sc_hd__mux2_1
Xfanout125 _3057_/A vssd1 vssd1 vccd1 vccd1 _3127_/A sky130_fd_sc_hd__buf_8
XANTENNA__2587__S _2589_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout114 _3112_/A vssd1 vssd1 vccd1 vccd1 _3101_/A sky130_fd_sc_hd__buf_8
X_3209_ _3333_/CLK _3209_/D vssd1 vssd1 vccd1 vccd1 _3209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold190 _3256_/Q vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2002__S0 _2045_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1890_ _1923_/A _2363_/A vssd1 vssd1 vccd1 vccd1 _2871_/C sky130_fd_sc_hd__nand2b_2
XFILLER_0_55_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3560_ _3576_/CLK _3560_/D _3054_/Y vssd1 vssd1 vccd1 vccd1 _3560_/Q sky130_fd_sc_hd__dfstp_1
X_2511_ hold82/A _2438_/B _2558_/C _3343_/Q _2509_/X vssd1 vssd1 vccd1 vccd1 _2511_/X
+ sky130_fd_sc_hd__o221a_1
X_3491_ _3602_/CLK _3491_/D _2985_/Y vssd1 vssd1 vccd1 vccd1 _3491_/Q sky130_fd_sc_hd__dfstp_1
X_2442_ _3512_/Q _2507_/C _2572_/A vssd1 vssd1 vccd1 vccd1 _2442_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2697__A1 _2406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2373_ _1825_/A _1793_/B _2370_/Y _3153_/Q vssd1 vssd1 vccd1 vccd1 _2373_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_75_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2544__S1 _1943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2870__S _2870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2709_ _2760_/A _2790_/B vssd1 vssd1 vccd1 vccd1 _2718_/S sky130_fd_sc_hd__or2_4
XANTENNA__2480__S0 _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2376__B1 _1769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2690__S _2697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2991_ _3049_/A vssd1 vssd1 vccd1 vccd1 _2991_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1942_ _3520_/Q _3519_/Q vssd1 vssd1 vccd1 vccd1 _1943_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_56_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1873_ _1845_/A _1845_/B _1837_/A vssd1 vssd1 vccd1 vccd1 _1873_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3612_ _3614_/CLK _3612_/D _3103_/Y vssd1 vssd1 vccd1 vccd1 _3612_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold904 _2379_/X vssd1 vssd1 vccd1 vccd1 hold904/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 _1872_/X vssd1 vssd1 vccd1 vccd1 _3530_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 _1884_/X vssd1 vssd1 vccd1 vccd1 _3524_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold915 _3569_/Q vssd1 vssd1 vccd1 vccd1 _1689_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3543_ _3573_/CLK _3543_/D _3037_/Y vssd1 vssd1 vccd1 vccd1 _3543_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3474_ _3533_/CLK _3474_/D _2968_/Y vssd1 vssd1 vccd1 vccd1 _3474_/Q sky130_fd_sc_hd__dfrtp_1
Xhold948 hold948/A vssd1 vssd1 vccd1 vccd1 _1742_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold959 _3556_/Q vssd1 vssd1 vccd1 vccd1 hold959/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_2_2__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2425_ _3634_/Q _2510_/A _2422_/X _2424_/X _2510_/B vssd1 vssd1 vccd1 vccd1 _2425_/X
+ sky130_fd_sc_hd__a221o_1
X_2356_ _3619_/Q _2356_/B vssd1 vssd1 vccd1 vccd1 _2363_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__2865__S _2870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2287_ hold35/A hold20/A vssd1 vssd1 vccd1 vccd1 _2510_/B sky130_fd_sc_hd__and2_4
XFILLER_0_59_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2775__S _2779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2597__A0 _2104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _2208_/Y _2210_/B _2210_/C vssd1 vssd1 vccd1 vccd1 _2210_/Y sky130_fd_sc_hd__nand3b_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _3431_/CLK _3190_/D vssd1 vssd1 vccd1 vccd1 _3190_/Q sky130_fd_sc_hd__dfxtp_1
X_2141_ _2139_/B _2140_/X _2143_/A _2119_/B vssd1 vssd1 vccd1 vccd1 _3497_/D sky130_fd_sc_hd__o2bb2a_1
X_2072_ _2058_/C _2069_/X _2070_/X _2090_/A _2067_/B vssd1 vssd1 vccd1 vccd1 _2072_/Y
+ sky130_fd_sc_hd__a2111oi_2
XFILLER_0_88_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2824__A1 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2974_ _3097_/A vssd1 vssd1 vccd1 vccd1 _2974_/Y sky130_fd_sc_hd__inv_2
X_1925_ _1929_/A _1932_/B vssd1 vssd1 vccd1 vccd1 _1934_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_6_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3332_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_16_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1856_ _1580_/Y _1837_/A _1853_/X _1855_/X vssd1 vssd1 vccd1 vccd1 _3538_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold701 _2600_/X vssd1 vssd1 vccd1 vccd1 _3146_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 _3157_/Q vssd1 vssd1 vccd1 vccd1 hold712/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1787_ _3554_/Q _2124_/B vssd1 vssd1 vccd1 vccd1 _1792_/B sky130_fd_sc_hd__xnor2_1
X_3526_ _3576_/CLK _3526_/D _3020_/Y vssd1 vssd1 vccd1 vccd1 _3526_/Q sky130_fd_sc_hd__dfrtp_1
Xhold745 _2882_/X vssd1 vssd1 vccd1 vccd1 _3412_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold734 _3191_/Q vssd1 vssd1 vccd1 vccd1 hold734/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 _2604_/X vssd1 vssd1 vccd1 vccd1 _3154_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout102_A hold45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold756 _3161_/Q vssd1 vssd1 vccd1 vccd1 hold756/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 _3579_/Q vssd1 vssd1 vccd1 vccd1 hold778/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 _2608_/X vssd1 vssd1 vccd1 vccd1 _3158_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3457_ _3594_/CLK _3457_/D _2951_/Y vssd1 vssd1 vccd1 vccd1 _3457_/Q sky130_fd_sc_hd__dfrtp_1
Xhold789 _1979_/X vssd1 vssd1 vccd1 vccd1 _3508_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3388_ _3433_/CLK _3388_/D vssd1 vssd1 vccd1 vccd1 _3388_/Q sky130_fd_sc_hd__dfxtp_1
X_2408_ _2165_/B _2421_/B hold63/A vssd1 vssd1 vccd1 vccd1 _2438_/B sky130_fd_sc_hd__o21ai_4
X_2339_ _3559_/Q _3558_/Q _3557_/Q _3556_/Q vssd1 vssd1 vccd1 vccd1 _2339_/X sky130_fd_sc_hd__or4_1
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2815__A1 _2104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold50 input3/X vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__buf_1
Xhold61 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__clkbuf_2
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2806__A1 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1710_ _3450_/Q _1865_/A vssd1 vssd1 vccd1 vccd1 _1710_/X sky130_fd_sc_hd__and2b_1
X_2690_ hold184/X _2802_/A1 _2697_/S vssd1 vssd1 vccd1 vccd1 _2690_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1641_ _2070_/A _2399_/A hold12/X vssd1 vssd1 vccd1 vccd1 _3621_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1572_ _1572_/A vssd1 vssd1 vccd1 vccd1 _1572_/Y sky130_fd_sc_hd__inv_2
X_3311_ _3320_/CLK _3311_/D vssd1 vssd1 vccd1 vccd1 _3311_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2742__A0 _2802_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ _3330_/CLK _3242_/D vssd1 vssd1 vccd1 vccd1 _3242_/Q sky130_fd_sc_hd__dfxtp_1
X_3173_ _3579_/CLK _3173_/D vssd1 vssd1 vccd1 vccd1 _3173_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2124_ _3498_/Q _2124_/B vssd1 vssd1 vccd1 vccd1 _2127_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__1613__A hold92/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2055_ hold804/X _2054_/Y _2055_/S vssd1 vssd1 vccd1 vccd1 _2055_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2957_ _3069_/A vssd1 vssd1 vccd1 vccd1 _2957_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2888_ _2072_/Y hold602/X _2890_/S vssd1 vssd1 vccd1 vccd1 _2888_/X sky130_fd_sc_hd__mux2_1
X_1908_ _1608_/A _3577_/Q _2577_/B _1908_/D vssd1 vssd1 vccd1 vccd1 _2162_/B sky130_fd_sc_hd__and4b_1
X_1839_ _1839_/A _1883_/A _3523_/Q vssd1 vssd1 vccd1 vccd1 _1879_/B sky130_fd_sc_hd__nand3_1
Xhold520 _3355_/Q vssd1 vssd1 vccd1 vccd1 hold520/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 _3425_/Q vssd1 vssd1 vccd1 vccd1 hold542/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 _2893_/X vssd1 vssd1 vccd1 vccd1 _3422_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 _2844_/X vssd1 vssd1 vccd1 vccd1 _3374_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold597 _2884_/X vssd1 vssd1 vccd1 vccd1 _3414_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 _3198_/Q vssd1 vssd1 vccd1 vccd1 hold586/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 _3176_/Q vssd1 vssd1 vccd1 vccd1 hold564/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 _2598_/X vssd1 vssd1 vccd1 vccd1 _3144_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3509_ _3509_/CLK _3509_/D _3003_/Y vssd1 vssd1 vccd1 vccd1 _3509_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2724__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput40 _3577_/Q vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_12
Xoutput51 _2453_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_12
Xoutput62 _2498_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_12
X_2811_ hold604/X _2358_/B _2819_/S vssd1 vssd1 vccd1 vccd1 _2811_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2742_ _2802_/A1 _2742_/A1 _2749_/S vssd1 vssd1 vccd1 vccd1 _2742_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2673_ hold303/X _2806_/A1 _2676_/S vssd1 vssd1 vccd1 vccd1 _2673_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2715__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1624_ _1624_/A _1624_/B hold18/X _1612_/B vssd1 vssd1 vccd1 vccd1 _1624_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_22_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1555_ _1767_/S vssd1 vssd1 vccd1 vccd1 _1689_/A sky130_fd_sc_hd__inv_2
X_3225_ _3333_/CLK _3225_/D vssd1 vssd1 vccd1 vccd1 _3225_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2479__C1 _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3156_ _3579_/CLK _3156_/D vssd1 vssd1 vccd1 vccd1 _3156_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2873__S _2880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2107_ _2064_/B _2088_/X _2091_/X _2064_/A _2067_/B vssd1 vssd1 vccd1 vccd1 _2107_/X
+ sky130_fd_sc_hd__a221o_1
X_3087_ _3090_/A vssd1 vssd1 vccd1 vccd1 _3087_/Y sky130_fd_sc_hd__inv_2
X_2038_ _3245_/Q _3317_/Q _3308_/Q _3299_/Q _2221_/B _2219_/A vssd1 vssd1 vccd1 vccd1
+ _2038_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2706__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold350 _2749_/X vssd1 vssd1 vccd1 vccd1 _3279_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 _3636_/Q vssd1 vssd1 vccd1 vccd1 _1888_/A sky130_fd_sc_hd__buf_1
Xhold372 _3318_/Q vssd1 vssd1 vccd1 vccd1 hold372/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 _3231_/Q vssd1 vssd1 vccd1 vccd1 hold394/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 _2803_/X vssd1 vssd1 vccd1 vccd1 _3327_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1050 _3440_/Q vssd1 vssd1 vccd1 vccd1 hold338/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2783__S hold38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3589_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_output63_A _2514_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1920__A1 _1912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3010_ _3110_/A vssd1 vssd1 vccd1 vccd1 _3010_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2693__S _2697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1610__B hold62/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2725_ _2806_/A1 hold376/X _2728_/S vssd1 vssd1 vccd1 vccd1 _2725_/X sky130_fd_sc_hd__mux2_1
X_2656_ _2708_/A _2729_/B vssd1 vssd1 vccd1 vccd1 _2800_/B sky130_fd_sc_hd__nand2_2
XANTENNA__2868__S _2870_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1607_ _1607_/A _1607_/B _1608_/A vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__and3_2
XFILLER_0_10_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2587_ hold435/X _2807_/A1 _2589_/S vssd1 vssd1 vccd1 vccd1 _2587_/X sky130_fd_sc_hd__mux2_1
Xfanout104 hold70/X vssd1 vssd1 vccd1 vccd1 _2806_/A1 sky130_fd_sc_hd__buf_4
Xfanout126 _3057_/A vssd1 vssd1 vccd1 vccd1 _3054_/A sky130_fd_sc_hd__buf_6
Xfanout115 _3112_/A vssd1 vssd1 vccd1 vccd1 _3110_/A sky130_fd_sc_hd__buf_8
X_3208_ _3330_/CLK _3208_/D vssd1 vssd1 vccd1 vccd1 _3208_/Q sky130_fd_sc_hd__dfxtp_1
X_3139_ _3438_/CLK _3139_/D vssd1 vssd1 vccd1 vccd1 _3139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2778__S _2779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 _2721_/X vssd1 vssd1 vccd1 vccd1 _3254_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold191 _2723_/X vssd1 vssd1 vccd1 vccd1 _3256_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2002__S1 _2045_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2018__S _2036_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2510_ _2510_/A _2510_/B vssd1 vssd1 vccd1 vccd1 _2559_/B sky130_fd_sc_hd__nor2_2
X_3490_ _3607_/CLK _3490_/D _2984_/Y vssd1 vssd1 vccd1 vccd1 _3490_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2441_ _3608_/Q _2435_/A _2439_/X _2440_/X _2420_/X vssd1 vssd1 vccd1 vccd1 _2441_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2372_ hold941/X _2379_/A _2372_/S vssd1 vssd1 vccd1 vccd1 _2372_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1767__S _1767_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2909__A0 _2355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2708_ _2708_/A _2729_/B vssd1 vssd1 vccd1 vccd1 _2790_/B sky130_fd_sc_hd__or2_2
XANTENNA__2480__S1 _1943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2639_ _2104_/B hold672/X _2643_/S vssd1 vssd1 vccd1 vccd1 _2639_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1991__S0 _2045_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2300__A1 hold70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2990_ _3049_/A vssd1 vssd1 vccd1 vccd1 _2990_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1941_ _1935_/Y _1935_/B _1941_/S vssd1 vssd1 vccd1 vccd1 _3511_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_83_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1872_ _1837_/A _1846_/Y _1871_/X _1871_/A _1836_/A vssd1 vssd1 vccd1 vccd1 _1872_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3611_ _3614_/CLK _3611_/D _3102_/Y vssd1 vssd1 vccd1 vccd1 _3611_/Q sky130_fd_sc_hd__dfrtp_1
Xhold927 _3527_/Q vssd1 vssd1 vccd1 vccd1 _1877_/A sky130_fd_sc_hd__clkbuf_2
Xhold916 _3528_/Q vssd1 vssd1 vccd1 vccd1 _1843_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_10_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3542_ _3573_/CLK _3542_/D _3036_/Y vssd1 vssd1 vccd1 vccd1 _3542_/Q sky130_fd_sc_hd__dfrtp_1
Xhold905 _2380_/X vssd1 vssd1 vccd1 vccd1 _3351_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3473_ _3567_/CLK _3473_/D _2967_/Y vssd1 vssd1 vccd1 vccd1 _3473_/Q sky130_fd_sc_hd__dfrtp_1
Xhold938 _3493_/Q vssd1 vssd1 vccd1 vccd1 _2129_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold949 _1819_/X vssd1 vssd1 vccd1 vccd1 hold949/X sky130_fd_sc_hd__dlygate4sd3_1
X_2424_ _2121_/A hold11/A _2423_/X _2572_/A vssd1 vssd1 vccd1 vccd1 _2424_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2355_ _3618_/Q _2355_/B vssd1 vssd1 vccd1 vccd1 _2363_/B sky130_fd_sc_hd__xnor2_1
X_2286_ hold19/X _2413_/B vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__nor2_2
XFILLER_0_79_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2791__S _2799_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3651__A _3655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2140_ _2119_/B _2139_/A _2000_/S vssd1 vssd1 vccd1 vccd1 _2140_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_56_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2071_ _2058_/C _2069_/X _2070_/X vssd1 vssd1 vccd1 vccd1 _2071_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_88_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2973_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2973_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1924_ _1924_/A _1924_/B _1929_/B vssd1 vssd1 vccd1 vccd1 _1935_/B sky130_fd_sc_hd__and3_1
XANTENNA__3098__A _3112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2588__A1 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1855_ _1855_/A _1858_/A vssd1 vssd1 vccd1 vccd1 _1855_/X sky130_fd_sc_hd__and2_1
XFILLER_0_71_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold702 _3183_/Q vssd1 vssd1 vccd1 vccd1 hold702/X sky130_fd_sc_hd__dlygate4sd3_1
X_1786_ _2121_/A _2065_/A _1785_/Y vssd1 vssd1 vccd1 vccd1 _2124_/B sky130_fd_sc_hd__o21ai_2
X_3525_ _3576_/CLK _3525_/D _3019_/Y vssd1 vssd1 vccd1 vccd1 _3525_/Q sky130_fd_sc_hd__dfrtp_1
Xhold724 _3430_/Q vssd1 vssd1 vccd1 vccd1 hold724/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 _2607_/X vssd1 vssd1 vccd1 vccd1 _3157_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 _3182_/Q vssd1 vssd1 vccd1 vccd1 hold746/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 _2647_/X vssd1 vssd1 vccd1 vccd1 _3191_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 _2611_/X vssd1 vssd1 vccd1 vccd1 _3161_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 _3362_/Q vssd1 vssd1 vccd1 vccd1 hold768/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold779 _2258_/X vssd1 vssd1 vccd1 vccd1 _3463_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3456_ _3594_/CLK _3456_/D _2950_/Y vssd1 vssd1 vccd1 vccd1 _3456_/Q sky130_fd_sc_hd__dfrtp_1
X_2407_ hold59/X hold98/A hold95/X vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__and3_1
X_3387_ _3434_/CLK _3387_/D vssd1 vssd1 vccd1 vccd1 _3387_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2876__S _2880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2338_ _2338_/A _2338_/B vssd1 vssd1 vccd1 vccd1 _2338_/Y sky130_fd_sc_hd__nor2_1
X_2269_ _2270_/B _2270_/C vssd1 vssd1 vccd1 vccd1 _2283_/B sky130_fd_sc_hd__and2_1
XFILLER_0_79_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2751__A1 _2801_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2786__S hold38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold93/X vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_45_wb_clk_i clkbuf_leaf_3_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3602_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3646__A _3655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1640_ _2063_/A _2400_/A hold12/X vssd1 vssd1 vccd1 vccd1 _3622_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1571_ _3610_/Q vssd1 vssd1 vccd1 vccd1 _1571_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3310_ _3320_/CLK _3310_/D vssd1 vssd1 vccd1 vccd1 _3310_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _3333_/CLK _3241_/D vssd1 vssd1 vccd1 vccd1 _3241_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2696__S _2697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3172_ _3516_/CLK _3172_/D vssd1 vssd1 vccd1 vccd1 _3172_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2123_ _2123_/A _2123_/B _2123_/C _2123_/D vssd1 vssd1 vccd1 vccd1 _2127_/A sky130_fd_sc_hd__and4_1
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2054_ _2144_/C _2319_/B _2053_/Y vssd1 vssd1 vccd1 vccd1 _2054_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2956_ _3069_/A vssd1 vssd1 vccd1 vccd1 _2956_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2887_ _2106_/X hold638/X _2890_/S vssd1 vssd1 vccd1 vccd1 _2887_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1907_ hold35/A _2421_/B vssd1 vssd1 vccd1 vccd1 _2574_/A sky130_fd_sc_hd__nand2_4
X_1838_ _1883_/A _3523_/Q vssd1 vssd1 vccd1 vccd1 _1838_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_32_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold510 _3354_/Q vssd1 vssd1 vccd1 vccd1 hold510/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2733__A1 _2803_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold543 _2896_/X vssd1 vssd1 vccd1 vccd1 _3425_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold521 _2823_/X vssd1 vssd1 vccd1 vccd1 _3355_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 _3169_/Q vssd1 vssd1 vccd1 vccd1 hold554/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 _3159_/Q vssd1 vssd1 vccd1 vccd1 hold532/X sky130_fd_sc_hd__dlygate4sd3_1
X_1769_ _1811_/S _1769_/B _2383_/B vssd1 vssd1 vccd1 vccd1 _1769_/X sky130_fd_sc_hd__or3_1
Xhold587 _2654_/X vssd1 vssd1 vccd1 vccd1 _3198_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 _2629_/X vssd1 vssd1 vccd1 vccd1 _3176_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 _3435_/Q vssd1 vssd1 vccd1 vccd1 hold576/X sky130_fd_sc_hd__dlygate4sd3_1
X_3508_ _3509_/CLK _3508_/D _3002_/Y vssd1 vssd1 vccd1 vccd1 _3508_/Q sky130_fd_sc_hd__dfrtp_1
Xhold598 _3415_/Q vssd1 vssd1 vccd1 vccd1 hold598/X sky130_fd_sc_hd__dlygate4sd3_1
X_3439_ _3550_/CLK _3439_/D _2933_/Y vssd1 vssd1 vccd1 vccd1 _3439_/Q sky130_fd_sc_hd__dfstp_2
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput52 _3649_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_12
Xoutput41 _2434_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_12
Xoutput63 _2514_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_12
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2660__A0 _2803_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2810_ _2891_/A _2810_/B vssd1 vssd1 vccd1 vccd1 _2819_/S sky130_fd_sc_hd__and2_4
X_2741_ _2801_/A1 hold226/X _2749_/S vssd1 vssd1 vccd1 vccd1 _2741_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2672_ hold449/X _2805_/A1 _2676_/S vssd1 vssd1 vccd1 vccd1 _2672_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1623_ hold92/A input3/X _1623_/C hold8/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__or4_1
X_3224_ _3333_/CLK _3224_/D vssd1 vssd1 vccd1 vccd1 _3224_/Q sky130_fd_sc_hd__dfxtp_1
.ends

