* NGSPICE file created from uart_macro_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

.subckt uart_macro_wrapper io_oeb[0] io_oeb[1] uart_irq uart_rx uart_tx vccd1 vssd1
+ wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3155_ _3423_/CLK _3155_/D vssd1 vssd1 vccd1 vccd1 _3155_/Q sky130_fd_sc_hd__dfxtp_1
X_2106_ _2106_/A _2106_/B vssd1 vssd1 vccd1 vccd1 _2107_/B sky130_fd_sc_hd__xnor2_1
X_3086_ _3105_/A vssd1 vssd1 vccd1 vccd1 _3086_/Y sky130_fd_sc_hd__inv_2
X_2037_ _2036_/X _2035_/X _2190_/A vssd1 vssd1 vccd1 vccd1 _2038_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_49_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2939_ _3128_/A vssd1 vssd1 vccd1 vccd1 _2939_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_72_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold362 _3219_/Q vssd1 vssd1 vccd1 vccd1 hold362/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 _3328_/Q vssd1 vssd1 vccd1 vccd1 hold351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold340 _2749_/X vssd1 vssd1 vccd1 vccd1 _3273_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 _2791_/X vssd1 vssd1 vccd1 vccd1 _3311_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold395 _2701_/X vssd1 vssd1 vccd1 vccd1 _3230_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 _3282_/Q vssd1 vssd1 vccd1 vccd1 hold384/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1040 _3642_/Q vssd1 vssd1 vccd1 vccd1 _1711_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2890__A0 _2109_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2642__A0 _2342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1684__A1 hold52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2881__A0 _2079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2633__A0 _2097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2724_ _2794_/B _2764_/A _2794_/A vssd1 vssd1 vccd1 vccd1 _2733_/S sky130_fd_sc_hd__or3b_4
XFILLER_0_14_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2655_ _2105_/B hold614/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2655_/X sky130_fd_sc_hd__mux2_1
X_1606_ _3065_/A vssd1 vssd1 vccd1 vccd1 _1606_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_10_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2586_ _2586_/A _2586_/B vssd1 vssd1 vccd1 vccd1 _2586_/Y sky130_fd_sc_hd__nor2_1
Xfanout127 _3131_/A vssd1 vssd1 vccd1 vccd1 _3128_/A sky130_fd_sc_hd__buf_8
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout116 _3044_/A vssd1 vssd1 vccd1 vccd1 _3073_/A sky130_fd_sc_hd__buf_8
Xfanout105 hold86/X vssd1 vssd1 vccd1 vccd1 _2809_/A1 sky130_fd_sc_hd__clkbuf_4
X_3207_ _3328_/CLK _3207_/D vssd1 vssd1 vccd1 vccd1 _3207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3138_ _3331_/CLK _3138_/D vssd1 vssd1 vccd1 vccd1 _3138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3069_ _3070_/A vssd1 vssd1 vccd1 vccd1 _3069_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2624__A0 _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1963__S _2045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold170 _2675_/X vssd1 vssd1 vccd1 vccd1 _3207_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _3216_/Q vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 _2726_/X vssd1 vssd1 vccd1 vccd1 _3252_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2863__A0 _2338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1666__A1 _2395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2615__A0 _2079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2034__S _2045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3654__A _3659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2440_ _3585_/Q hold67/A _2417_/B _3382_/Q vssd1 vssd1 vccd1 vccd1 _2440_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2371_ _3346_/Q _2366_/C _2370_/Y _2145_/D vssd1 vssd1 vccd1 vccd1 _2371_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_75_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2529__S0 _1911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2606__A0 _2075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout125_A _3131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2707_ _2807_/A1 hold227/X _2713_/S vssd1 vssd1 vccd1 vccd1 _2707_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2638_ _2075_/B hold762/X _2640_/S vssd1 vssd1 vccd1 vccd1 _2638_/X sky130_fd_sc_hd__mux2_1
X_2569_ _2511_/Y _2567_/Y _2581_/C _2511_/B _3454_/Q vssd1 vssd1 vccd1 vccd1 _2570_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_49_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1991__S1 _2222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2845__A0 _2342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1648__A1 hold49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2789__S _2793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1982__S1 _2193_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2836__A0 _2097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1639__A1 hold33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1940_ _1933_/Y _1933_/B _1940_/S vssd1 vssd1 vccd1 vccd1 _3515_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1871_ _1871_/A _1871_/B vssd1 vssd1 vccd1 vccd1 _1871_/X sky130_fd_sc_hd__or2_1
XFILLER_0_71_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3610_ _3610_/CLK _3610_/D _3101_/Y vssd1 vssd1 vccd1 vccd1 _3610_/Q sky130_fd_sc_hd__dfrtp_1
X_3541_ _3542_/CLK _3541_/D _3035_/Y vssd1 vssd1 vccd1 vccd1 _3541_/Q sky130_fd_sc_hd__dfrtp_1
Xhold917 _3468_/Q vssd1 vssd1 vccd1 vccd1 hold917/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold906 _2376_/X vssd1 vssd1 vccd1 vccd1 _3442_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold928 _2382_/X vssd1 vssd1 vccd1 vccd1 _3437_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3472_ _3579_/CLK _3472_/D _2966_/Y vssd1 vssd1 vccd1 vccd1 _3472_/Q sky130_fd_sc_hd__dfrtp_1
Xhold939 _2159_/X vssd1 vssd1 vccd1 vccd1 _3497_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2423_ _3606_/Q _2420_/Y _2421_/X _2422_/X vssd1 vssd1 vccd1 vccd1 _2423_/X sky130_fd_sc_hd__o211a_1
X_2354_ _1572_/Y _1931_/A _1891_/A _3343_/Q vssd1 vssd1 vccd1 vccd1 _2354_/X sky130_fd_sc_hd__a211o_1
X_2285_ _2285_/A _2285_/B vssd1 vssd1 vccd1 vccd1 _2285_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_74_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2070_ _2121_/A _3549_/Q _2089_/B _2069_/Y vssd1 vssd1 vccd1 vccd1 _2070_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_76_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2972_ _3065_/A vssd1 vssd1 vccd1 vccd1 _2972_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1923_ _1933_/A _1923_/B _1931_/B vssd1 vssd1 vccd1 vccd1 _1933_/B sky130_fd_sc_hd__and3b_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1854_ _1855_/B _1853_/X _1834_/A vssd1 vssd1 vccd1 vccd1 _1858_/A sky130_fd_sc_hd__o21ai_1
Xhold703 _2836_/X vssd1 vssd1 vccd1 vccd1 _3360_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1785_ _1797_/B _2124_/B vssd1 vssd1 vccd1 vccd1 _1791_/B sky130_fd_sc_hd__nand2_1
Xhold714 _3387_/Q vssd1 vssd1 vccd1 vccd1 hold714/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold725 _2839_/X vssd1 vssd1 vccd1 vccd1 _3363_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 _3367_/Q vssd1 vssd1 vccd1 vccd1 hold736/X sky130_fd_sc_hd__dlygate4sd3_1
X_3524_ _3526_/CLK _3524_/D _3018_/Y vssd1 vssd1 vccd1 vccd1 _3524_/Q sky130_fd_sc_hd__dfrtp_1
X_3455_ _3633_/CLK hold47/X _2949_/Y vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__dfrtp_1
Xhold758 _3177_/Q vssd1 vssd1 vccd1 vccd1 hold758/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 _2842_/X vssd1 vssd1 vccd1 vccd1 _3366_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold769 _2880_/X vssd1 vssd1 vccd1 vccd1 _3405_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2406_ _2407_/A hold19/A vssd1 vssd1 vccd1 vccd1 _2406_/X sky130_fd_sc_hd__and2_1
X_3386_ _3404_/CLK _3386_/D vssd1 vssd1 vccd1 vccd1 _3386_/Q sky130_fd_sc_hd__dfxtp_1
X_2337_ _2337_/A _2337_/B vssd1 vssd1 vccd1 vccd1 _2337_/Y sky130_fd_sc_hd__nor2_1
X_2268_ _2571_/A _3463_/Q _1593_/Y _3634_/Q _2267_/X vssd1 vssd1 vccd1 vccd1 _2268_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2892__S _2894_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2199_ _2196_/A _2189_/X _2196_/Y vssd1 vssd1 vccd1 vccd1 _3487_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2028__A1 _1985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2132__S _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__clkbuf_8
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__clkbuf_2
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__buf_2
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2019__A1 _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_14_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3488_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1570_ _1570_/A vssd1 vssd1 vccd1 vccd1 _1570_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2042__S _2053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _3493_/CLK _3240_/D vssd1 vssd1 vccd1 vccd1 _3240_/Q sky130_fd_sc_hd__dfxtp_1
X_3171_ _3582_/CLK _3171_/D vssd1 vssd1 vccd1 vccd1 _3171_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2122_ _3624_/Q _2134_/C vssd1 vssd1 vccd1 vccd1 _2123_/C sky130_fd_sc_hd__nand2_1
XANTENNA__1613__C _1625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2053_ hold828/X _2052_/X _2053_/S vssd1 vssd1 vccd1 vccd1 _2053_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2955_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2955_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2886_ _2096_/Y hold670/X _2894_/S vssd1 vssd1 vccd1 vccd1 _2886_/X sky130_fd_sc_hd__mux2_1
X_1906_ hold28/X hold19/X vssd1 vssd1 vccd1 vccd1 _2506_/S sky130_fd_sc_hd__and2_4
X_1837_ _1881_/A _1881_/B vssd1 vssd1 vccd1 vccd1 _1879_/B sky130_fd_sc_hd__or2_1
XFILLER_0_4_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold500 hold500/A vssd1 vssd1 vccd1 vccd1 _1928_/A sky130_fd_sc_hd__buf_1
Xhold511 _2333_/Y vssd1 vssd1 vccd1 vccd1 _3380_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 _3422_/Q vssd1 vssd1 vccd1 vccd1 hold544/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 _2827_/X vssd1 vssd1 vccd1 vccd1 _3352_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2887__S _2894_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold522 _3340_/Q vssd1 vssd1 vccd1 vccd1 hold522/X sky130_fd_sc_hd__dlygate4sd3_1
X_1768_ hold971/X _2383_/C _1767_/X vssd1 vssd1 vccd1 vccd1 _1768_/X sky130_fd_sc_hd__o21a_1
X_3507_ _3513_/CLK _3507_/D _3001_/Y vssd1 vssd1 vccd1 vccd1 _3507_/Q sky130_fd_sc_hd__dfrtp_1
X_1699_ _1700_/B _1700_/C _1698_/X vssd1 vssd1 vccd1 vccd1 _3578_/D sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold566 _3393_/Q vssd1 vssd1 vccd1 vccd1 hold566/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 _2898_/X vssd1 vssd1 vccd1 vccd1 _3421_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 _3149_/Q vssd1 vssd1 vccd1 vccd1 hold588/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 _2815_/X vssd1 vssd1 vccd1 vccd1 _3332_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold599 _2911_/X vssd1 vssd1 vccd1 vccd1 _3433_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3438_ _3551_/CLK _3438_/D _2932_/Y vssd1 vssd1 vccd1 vccd1 _3438_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _3369_/CLK _3369_/D vssd1 vssd1 vccd1 vccd1 _3369_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2497__A1 _3642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput42 _2570_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_12
Xoutput53 _3654_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_12
Xoutput64 _2535_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_12
XANTENNA__2098__A _2339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2032__S0 _2044_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3657__A _3659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2740_ _2810_/A1 hold325/X _2743_/S vssd1 vssd1 vccd1 vccd1 _2740_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2671_ _2812_/A1 hold327/X _2672_/S vssd1 vssd1 vccd1 vccd1 _2671_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1608__C _1907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1622_ _1559_/A _2395_/A _1623_/S vssd1 vssd1 vccd1 vccd1 _3639_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3223_ _3523_/CLK _3223_/D vssd1 vssd1 vccd1 vccd1 _3223_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1624__B input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3154_ _3582_/CLK _3154_/D vssd1 vssd1 vccd1 vccd1 _3154_/Q sky130_fd_sc_hd__dfxtp_1
X_3085_ _3124_/A vssd1 vssd1 vccd1 vccd1 _3085_/Y sky130_fd_sc_hd__inv_2
X_2105_ _2105_/A _2105_/B vssd1 vssd1 vccd1 vccd1 _2106_/B sky130_fd_sc_hd__xor2_1
X_2036_ hold171/X hold193/X hold187/X hold165/X _1590_/A _2222_/A vssd1 vssd1 vccd1
+ vccd1 _2036_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2938_ _3133_/A vssd1 vssd1 vccd1 vccd1 _2938_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2190__B _2222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2869_ hold534/X _2105_/B _2874_/S vssd1 vssd1 vccd1 vccd1 _2869_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold330 _2770_/X vssd1 vssd1 vccd1 vccd1 _3292_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 _2810_/X vssd1 vssd1 vccd1 vccd1 _3328_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 _3231_/Q vssd1 vssd1 vccd1 vccd1 hold341/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 _2689_/X vssd1 vssd1 vccd1 vccd1 _3219_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _3203_/Q vssd1 vssd1 vccd1 vccd1 hold374/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 _3240_/Q vssd1 vssd1 vccd1 vccd1 hold396/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 _2759_/X vssd1 vssd1 vccd1 vccd1 _3282_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2014__S0 _1590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1041 _3554_/Q vssd1 vssd1 vccd1 vccd1 _1806_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout68_A _2104_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1030 _3523_/Q vssd1 vssd1 vccd1 vccd1 _1905_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1052 _3348_/Q vssd1 vssd1 vccd1 vccd1 hold495/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2320__S _2320_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2556__A _3522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1610__D input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2723_ _2813_/A1 hold459/X _2723_/S vssd1 vssd1 vccd1 vccd1 _2723_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2654_ _2105_/A hold572/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2654_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1605_ _1808_/D vssd1 vssd1 vccd1 vccd1 _1605_/Y sky130_fd_sc_hd__inv_2
X_2585_ _2585_/A _2585_/B _2585_/C vssd1 vssd1 vccd1 vccd1 _2585_/X sky130_fd_sc_hd__and3_1
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout128 _3131_/A vssd1 vssd1 vccd1 vccd1 _3036_/A sky130_fd_sc_hd__buf_6
Xfanout117 _3044_/A vssd1 vssd1 vccd1 vccd1 _3070_/A sky130_fd_sc_hd__buf_4
Xfanout106 hold126/X vssd1 vssd1 vccd1 vccd1 _2808_/A1 sky130_fd_sc_hd__clkbuf_4
X_3206_ _3325_/CLK _3206_/D vssd1 vssd1 vccd1 vccd1 _3206_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2872__A1 _2075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3137_ _3328_/CLK _3137_/D vssd1 vssd1 vccd1 vccd1 _3137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3068_ _3070_/A vssd1 vssd1 vccd1 vccd1 _3068_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_54_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2019_ _3346_/Q _2017_/Y _2018_/Y vssd1 vssd1 vccd1 vccd1 _2019_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold171 _3243_/Q vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 _2665_/X vssd1 vssd1 vccd1 vccd1 _3198_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 _3315_/Q vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _2686_/X vssd1 vssd1 vccd1 vccd1 _3216_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2370_ _2370_/A vssd1 vssd1 vccd1 vccd1 _2370_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2529__S1 _2550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2706_ _2806_/A1 hold161/X _2713_/S vssd1 vssd1 vccd1 vccd1 _2706_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2790__A0 _2810_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2637_ _2079_/A hold750/X _2640_/S vssd1 vssd1 vccd1 vccd1 _2637_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout118_A _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2568_ hold67/A _2568_/B _2568_/C _2568_/D vssd1 vssd1 vccd1 vccd1 _2581_/C sky130_fd_sc_hd__and4_2
XFILLER_0_10_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2499_ _3372_/Q _3354_/Q _3363_/Q _3192_/Q _1943_/B _2550_/S1 vssd1 vssd1 vccd1 vccd1
+ _2499_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2781__A0 _2811_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_39_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3369_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2045__S _2045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1870_ _1835_/A _1847_/B _1869_/X _1845_/A _1560_/Y vssd1 vssd1 vccd1 vccd1 _1870_/X
+ sky130_fd_sc_hd__a32o_1
X_3540_ _3540_/CLK _3540_/D _3034_/Y vssd1 vssd1 vccd1 vccd1 _3540_/Q sky130_fd_sc_hd__dfrtp_1
Xhold918 _3535_/Q vssd1 vssd1 vccd1 vccd1 _1845_/A sky130_fd_sc_hd__buf_1
XANTENNA__2772__A0 _2812_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold907 _3576_/Q vssd1 vssd1 vccd1 vccd1 _1703_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3471_ _3579_/CLK _3471_/D _2965_/Y vssd1 vssd1 vccd1 vccd1 _3471_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold929 _3440_/Q vssd1 vssd1 vccd1 vccd1 _1815_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_2422_ _3607_/Q _2476_/B _2507_/C _3483_/Q vssd1 vssd1 vccd1 vccd1 _2422_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_19_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2353_ _1572_/Y _1931_/A _1928_/A _1573_/Y _2352_/X vssd1 vssd1 vccd1 vccd1 _2353_/X
+ sky130_fd_sc_hd__o221a_1
X_2284_ _2272_/A _2285_/B _2283_/Y vssd1 vssd1 vccd1 vccd1 _2284_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_79_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2827__A1 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1999_ hold392/X hold406/X hold410/X hold400/X _2044_/S0 _2044_/S1 vssd1 vssd1 vccd1
+ vccd1 _1999_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_15_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2818__A1 _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2429__S0 _1943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2506__A0 _2498_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2809__A1 _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2971_ _3065_/A vssd1 vssd1 vccd1 vccd1 _2971_/Y sky130_fd_sc_hd__inv_2
X_1922_ _2598_/C _1922_/B vssd1 vssd1 vccd1 vccd1 _1931_/B sky130_fd_sc_hd__nand2_4
X_1853_ _1853_/A _1859_/A _1859_/B vssd1 vssd1 vccd1 vccd1 _1853_/X sky130_fd_sc_hd__and3_1
XFILLER_0_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2745__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1784_ _1784_/A _1784_/B vssd1 vssd1 vccd1 vccd1 _2124_/B sky130_fd_sc_hd__nor2_1
Xhold715 _2860_/X vssd1 vssd1 vccd1 vccd1 _3387_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 _3386_/Q vssd1 vssd1 vccd1 vccd1 hold726/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold704 _3418_/Q vssd1 vssd1 vccd1 vccd1 hold704/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 _2843_/X vssd1 vssd1 vccd1 vccd1 _3367_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3523_ _3523_/CLK _3523_/D _3017_/Y vssd1 vssd1 vccd1 vccd1 _3523_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__1627__B _1668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3454_ _3637_/CLK hold3/X _2948_/Y vssd1 vssd1 vccd1 vccd1 _3454_/Q sky130_fd_sc_hd__dfrtp_2
Xhold759 _2639_/X vssd1 vssd1 vccd1 vccd1 _3177_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold748 _3159_/Q vssd1 vssd1 vccd1 vccd1 hold748/X sky130_fd_sc_hd__dlygate4sd3_1
X_2405_ _2071_/A _2571_/B _2511_/A vssd1 vssd1 vccd1 vccd1 _2405_/Y sky130_fd_sc_hd__a21oi_1
X_3385_ _3435_/CLK _3385_/D vssd1 vssd1 vccd1 vccd1 _3385_/Q sky130_fd_sc_hd__dfxtp_1
X_2336_ _3580_/Q _1889_/Y _3378_/Q vssd1 vssd1 vccd1 vccd1 _2337_/B sky130_fd_sc_hd__a21oi_1
X_2267_ hold38/A _2275_/A _3460_/Q _1563_/Y vssd1 vssd1 vccd1 vccd1 _2267_/X sky130_fd_sc_hd__a22o_1
X_2198_ _2222_/A _2196_/Y _2197_/Y _2196_/B vssd1 vssd1 vccd1 vccd1 _2198_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_47_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2736__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout98_A _2224_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__clkbuf_4
Xhold75 wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_85_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2019__A2 _2017_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2727__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _3423_/CLK _3170_/D vssd1 vssd1 vccd1 vccd1 _3170_/Q sky130_fd_sc_hd__dfxtp_1
X_2121_ _2121_/A _2134_/C vssd1 vssd1 vccd1 vccd1 _2123_/B sky130_fd_sc_hd__or2_1
X_2052_ hold820/X _2320_/S _2052_/S vssd1 vssd1 vccd1 vccd1 _2052_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2954_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2954_/Y sky130_fd_sc_hd__inv_2
X_2885_ _3526_/Q _2905_/B _2885_/C vssd1 vssd1 vccd1 vccd1 _2894_/S sky130_fd_sc_hd__or3_4
X_1905_ _1905_/A1 _2598_/C _1904_/Y vssd1 vssd1 vccd1 vccd1 _1905_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_44_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1836_ _1883_/A _3527_/Q vssd1 vssd1 vccd1 vccd1 _1881_/B sky130_fd_sc_hd__nand2_1
XANTENNA__2718__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold501 _3487_/Q vssd1 vssd1 vccd1 vccd1 hold501/X sky130_fd_sc_hd__dlygate4sd3_1
X_1767_ _1811_/A _1767_/B _1772_/B vssd1 vssd1 vccd1 vccd1 _1767_/X sky130_fd_sc_hd__or3_1
Xhold512 _3586_/Q vssd1 vssd1 vccd1 vccd1 hold512/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 _2899_/X vssd1 vssd1 vccd1 vccd1 _3422_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 _3395_/Q vssd1 vssd1 vccd1 vccd1 hold534/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 _2823_/X vssd1 vssd1 vccd1 vccd1 _3340_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3506_ _3623_/CLK _3506_/D _3000_/Y vssd1 vssd1 vccd1 vccd1 _3506_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1698_ _1700_/B _1700_/C _1700_/A vssd1 vssd1 vccd1 vccd1 _1698_/X sky130_fd_sc_hd__or3b_1
Xhold567 _2867_/X vssd1 vssd1 vccd1 vccd1 _3393_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 _3397_/Q vssd1 vssd1 vccd1 vccd1 hold556/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 _3389_/Q vssd1 vssd1 vccd1 vccd1 hold578/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold589 _2606_/X vssd1 vssd1 vccd1 vccd1 _3149_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3437_ _3580_/CLK _3437_/D _2931_/Y vssd1 vssd1 vccd1 vccd1 _3437_/Q sky130_fd_sc_hd__dfstp_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _3403_/CLK _3368_/D vssd1 vssd1 vccd1 vccd1 _3368_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2319_ _3624_/Q _2059_/A _2318_/X vssd1 vssd1 vccd1 vccd1 _2319_/X sky130_fd_sc_hd__o21ba_1
X_3299_ _3318_/CLK _3299_/D vssd1 vssd1 vccd1 vccd1 _3299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2709__A0 _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput43 _2573_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_12
Xoutput54 _3655_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_12
Xoutput65 _2548_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_12
XANTENNA__2032__S1 _2044_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2670_ _2811_/A1 hold374/X _2672_/S vssd1 vssd1 vccd1 vccd1 _2670_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2053__S _2053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1621_ _1558_/A _2396_/A _1623_/S vssd1 vssd1 vccd1 vccd1 _3640_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_1_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1624__C _1624_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3222_ _3612_/CLK _3222_/D vssd1 vssd1 vccd1 vccd1 _3222_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3153_ _3582_/CLK _3153_/D vssd1 vssd1 vccd1 vccd1 _3153_/Q sky130_fd_sc_hd__dfxtp_1
X_2104_ _2108_/A _2076_/C _2103_/X vssd1 vssd1 vccd1 vccd1 _2104_/X sky130_fd_sc_hd__o21a_2
XFILLER_0_27_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3084_ _3124_/A vssd1 vssd1 vccd1 vccd1 _3084_/Y sky130_fd_sc_hd__inv_2
X_2035_ _3288_/Q _3279_/Q _3270_/Q _3261_/Q _1590_/A _2222_/A vssd1 vssd1 vccd1 vccd1
+ _2035_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_57_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2937_ _3055_/A vssd1 vssd1 vccd1 vccd1 _2937_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2868_ hold538/X _2105_/A _2874_/S vssd1 vssd1 vccd1 vccd1 _2868_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2898__S _2904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2190__C _2224_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold320 _2780_/X vssd1 vssd1 vccd1 vccd1 _3301_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1819_ _1744_/A _1818_/X _1814_/X vssd1 vssd1 vccd1 vccd1 _1819_/X sky130_fd_sc_hd__o21a_1
X_2799_ hold424/X _2809_/A1 _2803_/S vssd1 vssd1 vccd1 vccd1 _2799_/X sky130_fd_sc_hd__mux2_1
Xhold331 _3274_/Q vssd1 vssd1 vccd1 vccd1 hold331/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1914__A1 _1911_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 _2702_/X vssd1 vssd1 vccd1 vccd1 _3231_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 _3222_/Q vssd1 vssd1 vccd1 vccd1 hold353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 _3320_/Q vssd1 vssd1 vccd1 vccd1 hold386/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 _2670_/X vssd1 vssd1 vccd1 vccd1 _3203_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 _3624_/Q vssd1 vssd1 vccd1 vccd1 hold364/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 _2712_/X vssd1 vssd1 vccd1 vccd1 _3240_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2014__S1 _2222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1020 _3477_/Q vssd1 vssd1 vccd1 vccd1 _2231_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 input18/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 _1905_/X vssd1 vssd1 vccd1 vccd1 _3523_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1053 _3349_/Q vssd1 vssd1 vccd1 vccd1 hold883/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1977__S _2052_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2722_ _2812_/A1 hold296/X _2723_/S vssd1 vssd1 vccd1 vccd1 _2722_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2653_ _2097_/A hold584/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2653_/X sky130_fd_sc_hd__mux2_1
X_1604_ _1824_/A vssd1 vssd1 vccd1 vccd1 _1604_/Y sky130_fd_sc_hd__inv_2
X_2584_ _2585_/A _2585_/B _2584_/C vssd1 vssd1 vccd1 vccd1 _2584_/X sky130_fd_sc_hd__and3_1
Xfanout129 _3089_/A vssd1 vssd1 vccd1 vccd1 _3131_/A sky130_fd_sc_hd__buf_4
XFILLER_0_1_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout118 _3089_/A vssd1 vssd1 vccd1 vccd1 _3044_/A sky130_fd_sc_hd__buf_4
Xfanout107 hold126/X vssd1 vssd1 vccd1 vccd1 _2397_/A sky130_fd_sc_hd__clkbuf_4
X_3205_ _3331_/CLK _3205_/D vssd1 vssd1 vccd1 vccd1 _3205_/Q sky130_fd_sc_hd__dfxtp_1
X_3136_ _3330_/CLK _3136_/D vssd1 vssd1 vccd1 vccd1 _3136_/Q sky130_fd_sc_hd__dfxtp_1
X_3067_ _3070_/A vssd1 vssd1 vccd1 vccd1 _3067_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2018_ _3509_/Q _3346_/Q vssd1 vssd1 vccd1 vccd1 _2018_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__1907__C_N _3581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold150 _3263_/Q vssd1 vssd1 vccd1 vccd1 hold150/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 _3234_/Q vssd1 vssd1 vccd1 vccd1 hold161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _2716_/X vssd1 vssd1 vccd1 vccd1 _3243_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 _2796_/X vssd1 vssd1 vccd1 vccd1 _3315_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _3324_/Q vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2303__A1 hold86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2506__S _2506_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold86_A hold86/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_9_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3325_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2705_ _2805_/A1 hold284/X _2713_/S vssd1 vssd1 vccd1 vccd1 _2705_/X sky130_fd_sc_hd__mux2_1
X_2636_ _2111_/B hold694/X _2640_/S vssd1 vssd1 vccd1 vccd1 _2636_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2567_ _2567_/A _2571_/B vssd1 vssd1 vccd1 vccd1 _2567_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_49_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2498_ hold88/A hold29/A _2496_/X _2497_/X vssd1 vssd1 vccd1 vccd1 _2498_/X sky130_fd_sc_hd__o22a_1
X_3119_ _3121_/A vssd1 vssd1 vccd1 vccd1 _3119_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1990__S _2045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold919 _1870_/X vssd1 vssd1 vccd1 vccd1 _3535_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold908 _1701_/B vssd1 vssd1 vccd1 vccd1 hold908/X sky130_fd_sc_hd__dlygate4sd3_1
X_3470_ _3579_/CLK _3470_/D _2964_/Y vssd1 vssd1 vccd1 vccd1 _3470_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2421_ _2413_/X _2414_/X _2417_/X _2441_/B _3595_/Q vssd1 vssd1 vccd1 vccd1 _2421_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__1958__S0 _2044_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2352_ _1575_/Y _1940_/S _2350_/X _2351_/X vssd1 vssd1 vccd1 vccd1 _2352_/X sky130_fd_sc_hd__a31o_1
X_2283_ _2285_/A _2283_/B vssd1 vssd1 vccd1 vccd1 _2283_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1998_ hold816/X _1997_/X _2053_/S vssd1 vssd1 vccd1 vccd1 _1998_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2763__A1 _2813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2619_ _3523_/Q _2630_/C _3524_/Q vssd1 vssd1 vccd1 vccd1 _2885_/C sky130_fd_sc_hd__or3b_2
X_3599_ _3614_/CLK _3599_/D _3090_/Y vssd1 vssd1 vccd1 vccd1 _3599_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2345__A2_N _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1985__S _1985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2429__S1 _1942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2690__A0 _2810_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2970_ _3105_/A vssd1 vssd1 vccd1 vccd1 _2970_/Y sky130_fd_sc_hd__inv_2
X_1921_ _1921_/A _2598_/C _1922_/B vssd1 vssd1 vccd1 vccd1 _1923_/B sky130_fd_sc_hd__or3_1
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1852_ _1859_/A _1859_/B vssd1 vssd1 vccd1 vccd1 _1852_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1783_ _1783_/A _2071_/A vssd1 vssd1 vccd1 vccd1 _1784_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_52_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold727 _2859_/X vssd1 vssd1 vccd1 vccd1 _3386_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold716 _3146_/Q vssd1 vssd1 vccd1 vccd1 hold716/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold705 _2894_/X vssd1 vssd1 vccd1 vccd1 _3418_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3522_ _3623_/CLK _3522_/D _3016_/Y vssd1 vssd1 vccd1 vccd1 _3522_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_52_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3453_ _3540_/CLK hold31/X _2947_/Y vssd1 vssd1 vccd1 vccd1 _3453_/Q sky130_fd_sc_hd__dfrtp_1
Xhold749 _2617_/X vssd1 vssd1 vccd1 vccd1 _3159_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 _3147_/Q vssd1 vssd1 vccd1 vccd1 hold738/X sky130_fd_sc_hd__dlygate4sd3_1
X_2404_ _2410_/A hold19/A hold28/A vssd1 vssd1 vccd1 vccd1 _2583_/B sky130_fd_sc_hd__o21ai_4
X_3384_ _3435_/CLK _3384_/D vssd1 vssd1 vccd1 vccd1 _3384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2335_ _2335_/A _2335_/B vssd1 vssd1 vccd1 vccd1 _2335_/Y sky130_fd_sc_hd__nor2_1
X_2266_ hold38/X _2275_/A _2273_/A _2571_/A _2265_/X vssd1 vssd1 vccd1 vccd1 _2269_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_46_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2197_ _2222_/A _2224_/B _2214_/A vssd1 vssd1 vccd1 vccd1 _2197_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold10 wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__clkbuf_4
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__buf_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__buf_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__buf_1
XANTENNA__2672__A0 _2813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3540_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2120_ _1588_/Y _2119_/X _1811_/A vssd1 vssd1 vccd1 vccd1 _2120_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2051_ _2051_/A vssd1 vssd1 vccd1 vccd1 _2320_/S sky130_fd_sc_hd__inv_2
X_2953_ _3128_/A vssd1 vssd1 vccd1 vccd1 _2953_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_72_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1904_ _1905_/A1 _2598_/C _1933_/A vssd1 vssd1 vccd1 vccd1 _1904_/Y sky130_fd_sc_hd__a21oi_1
X_2884_ _2339_/B hold672/X _2884_/S vssd1 vssd1 vccd1 vccd1 _2884_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1835_ _1835_/A vssd1 vssd1 vccd1 vccd1 _1855_/B sky130_fd_sc_hd__inv_2
Xhold502 _3490_/Q vssd1 vssd1 vccd1 vccd1 _2191_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1766_ _1763_/B _2383_/C _1765_/X vssd1 vssd1 vccd1 vccd1 _1766_/X sky130_fd_sc_hd__o21a_1
Xhold513 _2360_/Y vssd1 vssd1 vccd1 vccd1 _3342_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold535 _2869_/X vssd1 vssd1 vccd1 vccd1 _3395_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 _3392_/Q vssd1 vssd1 vccd1 vccd1 hold524/X sky130_fd_sc_hd__dlygate4sd3_1
X_3505_ _3551_/CLK _3505_/D _2999_/Y vssd1 vssd1 vccd1 vccd1 _3505_/Q sky130_fd_sc_hd__dfrtp_1
X_1697_ _1697_/A1 _1700_/C _1700_/A vssd1 vssd1 vccd1 vccd1 _1697_/X sky130_fd_sc_hd__o21a_1
Xhold546 _3350_/Q vssd1 vssd1 vccd1 vccd1 hold546/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 _3153_/Q vssd1 vssd1 vccd1 vccd1 hold568/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 _2871_/X vssd1 vssd1 vccd1 vccd1 _3397_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 _2862_/X vssd1 vssd1 vccd1 vccd1 _3389_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3436_ _3436_/CLK _3436_/D vssd1 vssd1 vccd1 vccd1 _3436_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _3526_/CLK _3367_/D vssd1 vssd1 vccd1 vccd1 _3367_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ _3627_/Q _2056_/A _2039_/Y vssd1 vssd1 vccd1 vccd1 _2318_/X sky130_fd_sc_hd__o21ba_1
X_3298_ _3316_/CLK _3298_/D vssd1 vssd1 vccd1 vccd1 _3298_/Q sky130_fd_sc_hd__dfxtp_1
X_2249_ _3474_/Q _3473_/Q _3472_/Q _3471_/Q vssd1 vssd1 vccd1 vccd1 _2250_/D sky130_fd_sc_hd__or4_1
XFILLER_0_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2654__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput55 _3656_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_12
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput66 _2562_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_12
Xoutput44 _2576_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_12
XANTENNA__2395__A _2395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2645__A0 _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1620__A1 _2397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1620_ _1770_/S _2397_/A _1623_/S vssd1 vssd1 vccd1 vccd1 _3641_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3221_ _3331_/CLK _3221_/D vssd1 vssd1 vccd1 vccd1 _3221_/Q sky130_fd_sc_hd__dfxtp_1
X_3152_ _3423_/CLK _3152_/D vssd1 vssd1 vccd1 vccd1 _3152_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2884__A0 _2339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1687__A1 _2397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2103_ _2056_/A _2090_/X _2102_/X _2076_/B vssd1 vssd1 vccd1 vccd1 _2103_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_27_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3083_ _3095_/A vssd1 vssd1 vccd1 vccd1 _3083_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2636__A0 _2111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2034_ _2032_/X _2033_/X _2045_/S vssd1 vssd1 vccd1 vccd1 _2034_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2936_ _3055_/A vssd1 vssd1 vccd1 vccd1 _2936_/Y sky130_fd_sc_hd__inv_2
X_2867_ hold566/X _2097_/A _2874_/S vssd1 vssd1 vccd1 vccd1 _2867_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1818_ _3555_/Q _1809_/B _1823_/A _3553_/Q vssd1 vssd1 vccd1 vccd1 _1818_/X sky130_fd_sc_hd__o211a_1
Xhold310 _2755_/X vssd1 vssd1 vccd1 vccd1 _3278_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2798_ hold185/X _2808_/A1 _2803_/S vssd1 vssd1 vccd1 vccd1 _2798_/X sky130_fd_sc_hd__mux2_1
Xhold332 _2750_/X vssd1 vssd1 vccd1 vccd1 _3274_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 _3283_/Q vssd1 vssd1 vccd1 vccd1 hold343/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 _3211_/Q vssd1 vssd1 vccd1 vccd1 hold321/X sky130_fd_sc_hd__dlygate4sd3_1
X_1749_ _1811_/A _1749_/B _1772_/B vssd1 vssd1 vccd1 vccd1 _1749_/X sky130_fd_sc_hd__or3_1
Xhold387 _2801_/X vssd1 vssd1 vccd1 vccd1 _3320_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1914__A2 _1911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold365 _1644_/X vssd1 vssd1 vccd1 vccd1 _3624_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 _3213_/Q vssd1 vssd1 vccd1 vccd1 hold376/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 _2692_/X vssd1 vssd1 vccd1 vccd1 _3222_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3419_ _3423_/CLK _3419_/D vssd1 vssd1 vccd1 vccd1 _3419_/Q sky130_fd_sc_hd__dfxtp_1
Xhold398 _3327_/Q vssd1 vssd1 vccd1 vccd1 hold398/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 _3464_/Q vssd1 vssd1 vccd1 vccd1 _2277_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1010 _2280_/Y vssd1 vssd1 vccd1 vccd1 _3463_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 _2241_/Y vssd1 vssd1 vccd1 vccd1 _3477_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1043 _1661_/C vssd1 vssd1 vccd1 vccd1 _1677_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold1054 _3606_/Q vssd1 vssd1 vccd1 vccd1 hold468/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2627__A0 _2075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1993__S _2045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3014__A _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2618__A0 _2339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2721_ _2811_/A1 hold355/X _2723_/S vssd1 vssd1 vccd1 vccd1 _2721_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2652_ _2342_/B hold706/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2652_/X sky130_fd_sc_hd__mux2_1
X_2583_ hold29/A _2583_/B _2583_/C vssd1 vssd1 vccd1 vccd1 _3659_/A sky130_fd_sc_hd__and3_4
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1603_ _1808_/B vssd1 vssd1 vccd1 vccd1 _1603_/Y sky130_fd_sc_hd__inv_2
Xfanout108 hold123/X vssd1 vssd1 vccd1 vccd1 _2807_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout119 _3121_/A vssd1 vssd1 vccd1 vccd1 _3055_/A sky130_fd_sc_hd__buf_6
X_3204_ _3330_/CLK _3204_/D vssd1 vssd1 vccd1 vccd1 _3204_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2857__A0 _2097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3135_ _3331_/CLK _3135_/D vssd1 vssd1 vccd1 vccd1 _3135_/Q sky130_fd_sc_hd__dfxtp_1
X_3066_ _3070_/A vssd1 vssd1 vccd1 vccd1 _3066_/Y sky130_fd_sc_hd__inv_2
X_2017_ _1985_/S _2012_/X _2016_/X vssd1 vssd1 vccd1 vccd1 _2017_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2919_ _3133_/A vssd1 vssd1 vccd1 vccd1 _2919_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_5_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold151 _2738_/X vssd1 vssd1 vccd1 vccd1 _3263_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold140 _3326_/Q vssd1 vssd1 vccd1 vccd1 hold140/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 _2706_/X vssd1 vssd1 vccd1 vccd1 _3234_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 input7/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _3270_/Q vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _2806_/X vssd1 vssd1 vccd1 vccd1 _3324_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2848__A0 _2104_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2612__S _2618_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2839__A0 _2111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2704_ _2794_/B _2784_/C _2794_/A vssd1 vssd1 vccd1 vccd1 _2713_/S sky130_fd_sc_hd__or3b_4
X_2635_ _2105_/B hold600/X _2640_/S vssd1 vssd1 vccd1 vccd1 _2635_/X sky130_fd_sc_hd__mux2_1
X_2566_ _2583_/B _2566_/B vssd1 vssd1 vccd1 vccd1 _2566_/X sky130_fd_sc_hd__and2_1
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2497_ _3642_/Q _2511_/A _2511_/B vssd1 vssd1 vccd1 vccd1 _2497_/X sky130_fd_sc_hd__a21o_1
X_3118_ _3121_/A vssd1 vssd1 vccd1 vccd1 _3118_/Y sky130_fd_sc_hd__inv_2
X_3049_ _3055_/A vssd1 vssd1 vccd1 vccd1 _3049_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_45_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_48_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3404_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout90 hold454/X vssd1 vssd1 vccd1 vccd1 _2794_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold909 _3587_/Q vssd1 vssd1 vccd1 vccd1 hold909/X sky130_fd_sc_hd__dlygate4sd3_1
X_2420_ _2584_/C vssd1 vssd1 vccd1 vccd1 _2420_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1958__S1 _2044_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2351_ _1573_/Y _1928_/A _2350_/B _2350_/A vssd1 vssd1 vccd1 vccd1 _2351_/X sky130_fd_sc_hd__a22o_1
X_2282_ _2273_/B _2283_/B _2281_/Y vssd1 vssd1 vccd1 vccd1 _3462_/D sky130_fd_sc_hd__o21a_1
XANTENNA__2517__S _2551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1997_ hold808/X _1996_/Y _2052_/S vssd1 vssd1 vccd1 vccd1 _1997_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout123_A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3598_ _3609_/CLK _3598_/D _3089_/Y vssd1 vssd1 vccd1 vccd1 _3598_/Q sky130_fd_sc_hd__dfrtp_1
X_2618_ _2339_/B hold610/X _2618_/S vssd1 vssd1 vccd1 vccd1 _2618_/X sky130_fd_sc_hd__mux2_1
X_2549_ _3409_/Q _3400_/Q _3391_/Q _3436_/Q _1911_/C _2550_/S1 vssd1 vssd1 vccd1 vccd1
+ _2549_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_65_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2398__A hold86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1920_ _1911_/C _1910_/Y _1917_/X vssd1 vssd1 vccd1 vccd1 _1920_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1851_ _1851_/A _1851_/B vssd1 vssd1 vccd1 vccd1 _1859_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3521_ _3623_/CLK _3521_/D _3015_/Y vssd1 vssd1 vccd1 vccd1 _3521_/Q sky130_fd_sc_hd__dfrtp_4
X_1782_ _3558_/Q _2126_/B vssd1 vssd1 vccd1 vccd1 _1791_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold717 _2603_/X vssd1 vssd1 vccd1 vccd1 _3146_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold728 _3414_/Q vssd1 vssd1 vccd1 vccd1 hold728/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold706 _3188_/Q vssd1 vssd1 vccd1 vccd1 hold706/X sky130_fd_sc_hd__dlygate4sd3_1
X_3452_ _3636_/CLK hold99/X _2946_/Y vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__dfrtp_1
Xhold739 _2604_/X vssd1 vssd1 vccd1 vccd1 _3147_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2403_ hold14/X _2403_/B vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__and2_1
X_3383_ _3523_/CLK _3383_/D vssd1 vssd1 vccd1 vccd1 _3383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2334_ _3504_/Q _1889_/Y _3379_/Q vssd1 vssd1 vccd1 vccd1 _2335_/B sky130_fd_sc_hd__a21oi_1
X_2265_ _3634_/Q _1593_/Y _3460_/Q _1563_/Y vssd1 vssd1 vccd1 vccd1 _2265_/X sky130_fd_sc_hd__o22a_1
X_2196_ _2196_/A _2196_/B vssd1 vssd1 vccd1 vccd1 _2196_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2681__A1 _2812_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2710__S _2713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2044__S0 _2044_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__clkbuf_4
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__buf_2
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__buf_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2035__S0 _1590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2050_ _1985_/S _2045_/X _2049_/X vssd1 vssd1 vccd1 vccd1 _2051_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2952_ _3128_/A vssd1 vssd1 vccd1 vccd1 _2952_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1903_ _2895_/C hold947/X _1933_/A vssd1 vssd1 vccd1 vccd1 _1903_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2883_ _2338_/B hold784/X _2884_/S vssd1 vssd1 vccd1 vccd1 _2883_/X sky130_fd_sc_hd__mux2_1
X_1834_ _1834_/A _1950_/B vssd1 vssd1 vccd1 vccd1 _1835_/A sky130_fd_sc_hd__and2_4
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1765_ _1811_/A _3561_/Q _1772_/B vssd1 vssd1 vccd1 vccd1 _1765_/X sky130_fd_sc_hd__or3_1
Xhold503 _2192_/X vssd1 vssd1 vccd1 vccd1 _3490_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 _3336_/Q vssd1 vssd1 vccd1 vccd1 hold536/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 _2866_/X vssd1 vssd1 vccd1 vccd1 _3392_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2530__S _2551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3504_ _3580_/CLK _3504_/D _2998_/Y vssd1 vssd1 vccd1 vccd1 _3504_/Q sky130_fd_sc_hd__dfrtp_1
Xhold514 _3588_/Q vssd1 vssd1 vccd1 vccd1 _2365_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 _2825_/X vssd1 vssd1 vccd1 vccd1 _3350_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3435_ _3435_/CLK _3435_/D vssd1 vssd1 vccd1 vccd1 _3435_/Q sky130_fd_sc_hd__dfxtp_1
X_1696_ _1701_/A _1701_/B vssd1 vssd1 vccd1 vccd1 _1700_/C sky130_fd_sc_hd__or2_2
Xhold569 _2611_/X vssd1 vssd1 vccd1 vccd1 _3153_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 _3428_/Q vssd1 vssd1 vccd1 vccd1 hold558/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3366_ _3369_/CLK _3366_/D vssd1 vssd1 vccd1 vccd1 _3366_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3297_ _3319_/CLK _3297_/D vssd1 vssd1 vccd1 vccd1 _3297_/Q sky130_fd_sc_hd__dfxtp_1
X_2317_ _2029_/Y _2315_/X _2316_/X vssd1 vssd1 vccd1 vccd1 _2323_/A sky130_fd_sc_hd__a21bo_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2248_ _3469_/Q _3468_/Q _3467_/Q _2247_/X _3475_/Q vssd1 vssd1 vccd1 vccd1 _2248_/X
+ sky130_fd_sc_hd__a41o_1
X_2179_ _2179_/A _3491_/Q _2661_/B vssd1 vssd1 vccd1 vccd1 _2804_/A sky130_fd_sc_hd__nand3_4
XANTENNA__2705__S _2713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1917__B1 _1911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput67 _2566_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_12
Xoutput56 _3657_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_12
Xoutput45 _2579_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_12
XFILLER_0_53_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2615__S _2618_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3220_ _3328_/CLK _3220_/D vssd1 vssd1 vccd1 vccd1 _3220_/Q sky130_fd_sc_hd__dfxtp_1
X_3151_ _3433_/CLK _3151_/D vssd1 vssd1 vccd1 vccd1 _3151_/Q sky130_fd_sc_hd__dfxtp_1
X_2102_ _2071_/A _3549_/Q _2089_/B _2062_/Y _2056_/B vssd1 vssd1 vccd1 vccd1 _2102_/X
+ sky130_fd_sc_hd__a311o_1
X_3082_ _3133_/A vssd1 vssd1 vccd1 vccd1 _3082_/Y sky130_fd_sc_hd__inv_2
X_2033_ hold181/X hold169/X hold159/X hold183/X _2044_/S0 _2044_/S1 vssd1 vssd1 vccd1
+ vccd1 _2033_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2935_ _3055_/A vssd1 vssd1 vccd1 vccd1 _2935_/Y sky130_fd_sc_hd__inv_2
X_2866_ hold524/X _2342_/B _2874_/S vssd1 vssd1 vccd1 vccd1 _2866_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1817_ _1817_/A _1817_/B vssd1 vssd1 vccd1 vccd1 _1823_/A sky130_fd_sc_hd__nor2_1
X_2797_ hold233/X _2807_/A1 _2803_/S vssd1 vssd1 vccd1 vccd1 _2797_/X sky130_fd_sc_hd__mux2_1
Xhold300 _3285_/Q vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold311 _3229_/Q vssd1 vssd1 vccd1 vccd1 hold311/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 _2760_/X vssd1 vssd1 vccd1 vccd1 _3283_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 _3266_/Q vssd1 vssd1 vccd1 vccd1 hold333/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold322 _2679_/X vssd1 vssd1 vccd1 vccd1 _3211_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1748_ hold925/X _2383_/C _1747_/X vssd1 vssd1 vccd1 vccd1 _1748_/X sky130_fd_sc_hd__o21a_1
Xhold366 _3286_/Q vssd1 vssd1 vccd1 vccd1 hold366/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 _3248_/Q vssd1 vssd1 vccd1 vccd1 hold355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 _2681_/X vssd1 vssd1 vccd1 vccd1 _3213_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1679_ hold19/X _2415_/A vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__nand2_1
X_3418_ _3427_/CLK _3418_/D vssd1 vssd1 vccd1 vccd1 _3418_/Q sky130_fd_sc_hd__dfxtp_1
Xhold399 _2809_/X vssd1 vssd1 vccd1 vccd1 _3327_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 _3291_/Q vssd1 vssd1 vccd1 vccd1 hold388/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1000 _3480_/Q vssd1 vssd1 vccd1 vccd1 _2261_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3349_ _3580_/CLK _3349_/D _2924_/Y vssd1 vssd1 vccd1 vccd1 _3349_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1033 _2278_/X vssd1 vssd1 vccd1 vccd1 _3464_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1011 _3462_/Q vssd1 vssd1 vccd1 vccd1 _2273_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1022 _3527_/Q vssd1 vssd1 vccd1 vccd1 _1885_/S sky130_fd_sc_hd__dlygate4sd3_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1044 _2415_/A vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1055 _3641_/Q vssd1 vssd1 vccd1 vccd1 hold208/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2866__A1 _2342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2720_ _2810_/A1 hold305/X _2723_/S vssd1 vssd1 vccd1 vccd1 _2720_/X sky130_fd_sc_hd__mux2_1
X_2651_ _2824_/B _2905_/B _2905_/C vssd1 vssd1 vccd1 vccd1 _2660_/S sky130_fd_sc_hd__nand3_4
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1602_ _1808_/A vssd1 vssd1 vccd1 vccd1 _1602_/Y sky130_fd_sc_hd__inv_2
X_2582_ _3459_/Q hold29/A _2583_/B _2583_/C vssd1 vssd1 vccd1 vccd1 _2582_/X sky130_fd_sc_hd__o211a_1
Xfanout109 hold123/X vssd1 vssd1 vccd1 vccd1 _2396_/A sky130_fd_sc_hd__clkbuf_4
X_3203_ _3331_/CLK _3203_/D vssd1 vssd1 vccd1 vccd1 _3203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3134_ _3493_/CLK _3134_/D vssd1 vssd1 vccd1 vccd1 _3134_/Q sky130_fd_sc_hd__dfxtp_1
X_3065_ _3065_/A vssd1 vssd1 vccd1 vccd1 _3065_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_54_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2016_ _1985_/S _2016_/B vssd1 vssd1 vccd1 vccd1 _2016_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2918_ _3105_/A vssd1 vssd1 vccd1 vccd1 _2918_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2793__A0 _2813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2849_ _2111_/B hold674/X _2853_/S vssd1 vssd1 vccd1 vccd1 _2849_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_13_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold141 _2808_/X vssd1 vssd1 vccd1 vccd1 _3326_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 _3218_/Q vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 _3225_/Q vssd1 vssd1 vccd1 vccd1 hold152/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 _2746_/X vssd1 vssd1 vccd1 vccd1 _3270_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _3317_/Q vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 _3308_/Q vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 input7/X vssd1 vssd1 vccd1 vccd1 _1659_/A sky130_fd_sc_hd__buf_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2583__B _2583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2775__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2703_ _2813_/A1 hold440/X _2703_/S vssd1 vssd1 vccd1 vccd1 _2703_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2634_ _2105_/A hold642/X _2640_/S vssd1 vssd1 vccd1 vccd1 _2634_/X sky130_fd_sc_hd__mux2_1
X_2565_ _3453_/Q _2511_/B _2568_/D _2564_/X vssd1 vssd1 vccd1 vccd1 _2566_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_49_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2496_ _3628_/Q hold7/A _2492_/X _2495_/X vssd1 vssd1 vccd1 vccd1 _2496_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_4_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3117_ _3121_/A vssd1 vssd1 vccd1 vccd1 _3117_/Y sky130_fd_sc_hd__inv_2
X_3048_ _3070_/A vssd1 vssd1 vccd1 vccd1 _3048_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2713__S _2713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2766__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2623__S _2629_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout91 hold259/X vssd1 vssd1 vccd1 vccd1 _2794_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3610_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2350_ _2350_/A _2350_/B vssd1 vssd1 vccd1 vccd1 _2350_/X sky130_fd_sc_hd__or2_1
X_2281_ _2273_/B _2283_/B _2285_/A vssd1 vssd1 vccd1 vccd1 _2281_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__1732__B2 _1595_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2748__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2533__S _2551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1996_ _1996_/A vssd1 vssd1 vccd1 vccd1 _1996_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_51_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3597_ _3633_/CLK _3597_/D _3088_/Y vssd1 vssd1 vccd1 vccd1 _3597_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2617_ _2338_/B hold748/X _2618_/S vssd1 vssd1 vccd1 vccd1 _2617_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2548_ _2583_/B _2540_/X _2547_/X _2506_/S vssd1 vssd1 vccd1 vccd1 _2548_/X sky130_fd_sc_hd__a22o_1
X_2479_ _3486_/Q _2507_/C _2476_/Y _2478_/X _2508_/A vssd1 vssd1 vccd1 vccd1 _2479_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__2708__S _2713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2739__A0 _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2911__A0 _2079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2618__S _2618_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1850_ _1850_/A vssd1 vssd1 vccd1 vccd1 _1851_/B sky130_fd_sc_hd__inv_2
XFILLER_0_21_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1781_ _3624_/Q _2056_/A _1780_/Y vssd1 vssd1 vccd1 vccd1 _2126_/B sky130_fd_sc_hd__o21ai_2
X_3520_ _3623_/CLK _3520_/D _3014_/Y vssd1 vssd1 vccd1 vccd1 _3520_/Q sky130_fd_sc_hd__dfrtp_1
Xhold718 _3388_/Q vssd1 vssd1 vccd1 vccd1 hold718/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold707 _2652_/X vssd1 vssd1 vccd1 vccd1 _3188_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3451_ _3540_/CLK hold63/X _2945_/Y vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__dfrtp_1
Xhold729 _2890_/X vssd1 vssd1 vccd1 vccd1 _3414_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3382_ _3633_/CLK _3382_/D _2930_/Y vssd1 vssd1 vccd1 vccd1 _3382_/Q sky130_fd_sc_hd__dfrtp_1
X_2402_ hold49/X _2403_/B vssd1 vssd1 vccd1 vccd1 _3592_/D sky130_fd_sc_hd__and2_1
X_2333_ _2333_/A _2333_/B vssd1 vssd1 vccd1 vccd1 _2333_/Y sky130_fd_sc_hd__nor2_1
X_2264_ hold23/X _2272_/A vssd1 vssd1 vccd1 vccd1 _2269_/B sky130_fd_sc_hd__xnor2_1
X_2195_ _2189_/X _2244_/B _2190_/A _2196_/B vssd1 vssd1 vccd1 vccd1 _2195_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1668__A _1668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2197__A1 _2222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1979_ _3257_/Q hold445/X hold426/X _3230_/Q _2224_/B _2193_/A1 vssd1 vssd1 vccd1
+ vccd1 _1979_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_70_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2044__S1 _2044_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 input3/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__buf_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3123__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2901__S _2904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2035__S1 _2222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2951_ _3128_/A vssd1 vssd1 vccd1 vccd1 _2951_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_69_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1902_ _1902_/A _1902_/B vssd1 vssd1 vccd1 vccd1 _1902_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_32_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3551_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2882_ _2075_/B hold560/X _2884_/S vssd1 vssd1 vccd1 vccd1 _2882_/X sky130_fd_sc_hd__mux2_1
X_1833_ _3544_/Q hold888/X _1833_/S vssd1 vssd1 vccd1 vccd1 _1833_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2811__S _2813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1764_ _1761_/B _1745_/Y _1763_/X vssd1 vssd1 vccd1 vccd1 _1764_/X sky130_fd_sc_hd__o21a_1
Xhold504 _3489_/Q vssd1 vssd1 vccd1 vccd1 _2190_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold526 _3351_/Q vssd1 vssd1 vccd1 vccd1 hold526/X sky130_fd_sc_hd__dlygate4sd3_1
X_3503_ _3551_/CLK _3503_/D _2997_/Y vssd1 vssd1 vccd1 vccd1 _3503_/Q sky130_fd_sc_hd__dfrtp_1
Xhold515 _2365_/Y vssd1 vssd1 vccd1 vccd1 _3341_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 _3353_/Q vssd1 vssd1 vccd1 vccd1 hold548/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 _2819_/X vssd1 vssd1 vccd1 vccd1 _3336_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1695_ _1703_/A _1703_/B vssd1 vssd1 vccd1 vccd1 _1701_/B sky130_fd_sc_hd__or2_1
Xhold559 _2906_/X vssd1 vssd1 vccd1 vccd1 _3428_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3434_ _3436_/CLK _3434_/D vssd1 vssd1 vccd1 vccd1 _3434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _3416_/CLK _3365_/D vssd1 vssd1 vccd1 vccd1 _3365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _3316_/CLK _3296_/D vssd1 vssd1 vccd1 vccd1 _3296_/Q sky130_fd_sc_hd__dfxtp_1
X_2316_ _3627_/Q _3626_/Q _1784_/B _2029_/Y _2315_/X vssd1 vssd1 vccd1 vccd1 _2316_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2247_ _3474_/Q _3473_/Q _3472_/Q _3471_/Q vssd1 vssd1 vccd1 vccd1 _2247_/X sky130_fd_sc_hd__and4_1
XFILLER_0_79_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2178_ _3491_/Q _2661_/B _2179_/A vssd1 vssd1 vccd1 vccd1 _2178_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_67_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2590__A1 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput57 _3658_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_12
Xoutput46 _2580_/Y vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_12
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3150_ _3435_/CLK _3150_/D vssd1 vssd1 vccd1 vccd1 _3150_/Q sky130_fd_sc_hd__dfxtp_1
X_3081_ _3133_/A vssd1 vssd1 vccd1 vccd1 _3081_/Y sky130_fd_sc_hd__inv_2
X_2101_ _2108_/A _2073_/X _2100_/Y _2076_/B vssd1 vssd1 vccd1 vccd1 _2101_/X sky130_fd_sc_hd__o211a_1
X_2032_ hold191/X hold202/X hold161/X hold152/X _2044_/S0 _2044_/S1 vssd1 vssd1 vccd1
+ vccd1 _2032_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2806__S _2813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2934_ _3055_/A vssd1 vssd1 vccd1 vccd1 _2934_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2865_ _2895_/C _2875_/B vssd1 vssd1 vccd1 vccd1 _2874_/S sky130_fd_sc_hd__nor2_4
X_1816_ _1745_/B _1813_/Y _1814_/X _1815_/X vssd1 vssd1 vccd1 vccd1 _1816_/X sky130_fd_sc_hd__o22a_1
Xhold301 _2762_/X vssd1 vssd1 vccd1 vccd1 _3285_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2796_ hold193/X _2806_/A1 _2803_/S vssd1 vssd1 vccd1 vccd1 _2796_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold334 _2741_/X vssd1 vssd1 vccd1 vccd1 _3266_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 _3202_/Q vssd1 vssd1 vccd1 vccd1 hold323/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 _2700_/X vssd1 vssd1 vccd1 vccd1 _3229_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1747_ _1811_/A _3570_/Q _1772_/B vssd1 vssd1 vccd1 vccd1 _1747_/X sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold378 _3304_/Q vssd1 vssd1 vccd1 vccd1 hold378/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 _2763_/X vssd1 vssd1 vccd1 vccd1 _3286_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 _2721_/X vssd1 vssd1 vccd1 vccd1 _3248_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold345 _3141_/Q vssd1 vssd1 vccd1 vccd1 hold345/X sky130_fd_sc_hd__dlygate4sd3_1
X_1678_ hold19/A _2415_/A vssd1 vssd1 vccd1 vccd1 _1678_/X sky130_fd_sc_hd__and2_1
X_3417_ _3583_/CLK _3417_/D vssd1 vssd1 vccd1 vccd1 _3417_/Q sky130_fd_sc_hd__dfxtp_1
Xhold389 _2769_/X vssd1 vssd1 vccd1 vccd1 _3291_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3348_ _3580_/CLK _3348_/D _2923_/Y vssd1 vssd1 vccd1 vccd1 _3348_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 _2235_/X vssd1 vssd1 vccd1 vccd1 _2236_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1023 _3502_/Q vssd1 vssd1 vccd1 vccd1 _2134_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1012 _3496_/Q vssd1 vssd1 vccd1 vccd1 _2160_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1045 _2396_/X vssd1 vssd1 vccd1 vccd1 _3586_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3279_ _3319_/CLK _3279_/D vssd1 vssd1 vccd1 vccd1 _3279_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1034 _3582_/Q vssd1 vssd1 vccd1 vccd1 hold478/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1056 _3347_/Q vssd1 vssd1 vccd1 vccd1 hold1056/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold890 _3344_/Q vssd1 vssd1 vccd1 vccd1 _1956_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__2626__S _2629_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2650_ _2339_/B hold664/X _2650_/S vssd1 vssd1 vccd1 vccd1 _2650_/X sky130_fd_sc_hd__mux2_1
X_1601_ _1956_/B vssd1 vssd1 vccd1 vccd1 _1601_/Y sky130_fd_sc_hd__inv_2
X_2581_ hold96/A hold7/A _2581_/C vssd1 vssd1 vccd1 vccd1 _2583_/C sky130_fd_sc_hd__and3_1
XANTENNA__1988__S0 _2044_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2306__A1 _2395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3202_ _3328_/CLK _3202_/D vssd1 vssd1 vccd1 vccd1 _3202_/Q sky130_fd_sc_hd__dfxtp_1
X_3133_ _3133_/A vssd1 vssd1 vccd1 vccd1 _3133_/Y sky130_fd_sc_hd__inv_2
X_3064_ _3131_/A vssd1 vssd1 vccd1 vccd1 _3064_/Y sky130_fd_sc_hd__inv_2
X_2015_ _2014_/X _2013_/X _2045_/S vssd1 vssd1 vccd1 vccd1 _2016_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_45_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2917_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2917_/Y sky130_fd_sc_hd__inv_2
X_2848_ _2104_/X hold708/X _2853_/S vssd1 vssd1 vccd1 vccd1 _2848_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2779_ _2809_/A1 hold414/X _2783_/S vssd1 vssd1 vccd1 vccd1 _2779_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold120 input27/X vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__clkbuf_2
Xhold142 _3209_/Q vssd1 vssd1 vccd1 vccd1 hold142/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 _2688_/X vssd1 vssd1 vccd1 vccd1 _3218_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 _2696_/X vssd1 vssd1 vccd1 vccd1 _3225_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1979__S0 _2224_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold175 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 input20/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _2788_/X vssd1 vssd1 vccd1 vccd1 _3308_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 _2798_/X vssd1 vssd1 vccd1 vccd1 _3317_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 _1677_/B vssd1 vssd1 vccd1 vccd1 _1661_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3131__A _3131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2702_ _2812_/A1 hold341/X _2703_/S vssd1 vssd1 vccd1 vccd1 _2702_/X sky130_fd_sc_hd__mux2_1
X_2633_ _2097_/A hold650/X _2640_/S vssd1 vssd1 vccd1 vccd1 _2633_/X sky130_fd_sc_hd__mux2_1
X_2564_ _3605_/Q _2568_/B _2417_/B _3381_/Q _2563_/X vssd1 vssd1 vccd1 vccd1 _2564_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1943__B _1943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2495_ _3619_/Q _1645_/Y _2493_/Y _2494_/X _2571_/B vssd1 vssd1 vccd1 vccd1 _2495_/X
+ sky130_fd_sc_hd__a221o_1
X_3116_ _3121_/A vssd1 vssd1 vccd1 vccd1 _3116_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3047_ _3070_/A vssd1 vssd1 vccd1 vccd1 _3047_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_81_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3126__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2904__S _2904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2757__A1 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout70 _2109_/X vssd1 vssd1 vccd1 vccd1 _2111_/B sky130_fd_sc_hd__buf_4
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout81 hold364/X vssd1 vssd1 vccd1 vccd1 _2121_/A sky130_fd_sc_hd__buf_4
Xfanout92 _2191_/A vssd1 vssd1 vccd1 vccd1 _1985_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2280_ _2285_/A _2280_/B _2280_/C vssd1 vssd1 vccd1 vccd1 _2280_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_19_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2693__A0 _2813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1995_ _1985_/S _1990_/X _1994_/X vssd1 vssd1 vccd1 vccd1 _1996_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_70_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2616_ _2075_/B hold648/X _2618_/S vssd1 vssd1 vccd1 vccd1 _2616_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout109_A hold123/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3596_ _3609_/CLK _3596_/D _3087_/Y vssd1 vssd1 vccd1 vccd1 _3596_/Q sky130_fd_sc_hd__dfrtp_1
X_2547_ _2546_/X _2543_/X _3522_/Q vssd1 vssd1 vccd1 vccd1 _2547_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2478_ _3587_/Q hold67/A _2508_/B _2477_/X vssd1 vssd1 vccd1 vccd1 _2478_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_76_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2531__S0 _2554_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2427__B1 _2583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2634__S _2640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1650__A1 hold52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1780_ _3625_/Q _3624_/Q _3626_/Q vssd1 vssd1 vccd1 vccd1 _1780_/Y sky130_fd_sc_hd__o21ai_1
Xhold708 _3371_/Q vssd1 vssd1 vccd1 vccd1 hold708/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold719 _2861_/X vssd1 vssd1 vccd1 vccd1 _3388_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3450_ _3499_/CLK _3450_/D _2944_/Y vssd1 vssd1 vccd1 vccd1 _3450_/Q sky130_fd_sc_hd__dfrtp_1
X_3381_ _3540_/CLK _3381_/D _2929_/Y vssd1 vssd1 vccd1 vccd1 _3381_/Q sky130_fd_sc_hd__dfrtp_1
X_2401_ hold44/X _2403_/B vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__and2_1
X_2332_ _1891_/A _1889_/Y _3380_/Q vssd1 vssd1 vccd1 vccd1 _2333_/B sky130_fd_sc_hd__a21oi_1
X_2263_ _2263_/A _2263_/B vssd1 vssd1 vccd1 vccd1 _2269_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__2809__S _2813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2666__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2194_ _2194_/A _2194_/B vssd1 vssd1 vccd1 vccd1 _2244_/B sky130_fd_sc_hd__or2_1
XANTENNA__1641__A1 _2397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2197__A2 _2224_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1978_ hold810/X _1977_/X _2053_/S vssd1 vssd1 vccd1 vccd1 _1978_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3579_ _3579_/CLK _3579_/D _3073_/Y vssd1 vssd1 vccd1 vccd1 _3579_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold13 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3328_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2657__A0 _2079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold57 input3/X vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__buf_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2454__S _3522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2629__S _2629_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2648__A0 _2075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2950_ _3128_/A vssd1 vssd1 vccd1 vccd1 _2950_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2881_ _2079_/A hold782/X _2884_/S vssd1 vssd1 vccd1 vccd1 _2881_/X sky130_fd_sc_hd__mux2_1
X_1901_ _1902_/A _1902_/B vssd1 vssd1 vccd1 vccd1 _2895_/C sky130_fd_sc_hd__or2_4
XFILLER_0_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1623__A1 _2585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1832_ hold877/X _3544_/Q _1833_/S vssd1 vssd1 vccd1 vccd1 _1832_/X sky130_fd_sc_hd__mux2_1
X_1763_ _1811_/A _1763_/B _1772_/B vssd1 vssd1 vccd1 vccd1 _1763_/X sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold505 _2195_/X vssd1 vssd1 vccd1 vccd1 _3489_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 _2826_/X vssd1 vssd1 vccd1 vccd1 _3351_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1694_ _1705_/A _1705_/B vssd1 vssd1 vccd1 vccd1 _1703_/B sky130_fd_sc_hd__or2_1
Xhold516 _3398_/Q vssd1 vssd1 vccd1 vccd1 hold516/X sky130_fd_sc_hd__dlygate4sd3_1
X_3502_ _3551_/CLK _3502_/D _2996_/Y vssd1 vssd1 vccd1 vccd1 _3502_/Q sky130_fd_sc_hd__dfrtp_1
Xhold549 _2828_/X vssd1 vssd1 vccd1 vccd1 _3353_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3433_ _3433_/CLK _3433_/D vssd1 vssd1 vccd1 vccd1 _3433_/Q sky130_fd_sc_hd__dfxtp_1
Xhold538 _3394_/Q vssd1 vssd1 vccd1 vccd1 hold538/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _3416_/CLK _3364_/D vssd1 vssd1 vccd1 vccd1 _3364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3295_ _3483_/CLK _3295_/D vssd1 vssd1 vccd1 vccd1 _3295_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2315_ _3627_/Q _3626_/Q _2017_/Y vssd1 vssd1 vccd1 vccd1 _2315_/X sky130_fd_sc_hd__o21ba_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2639__A0 _2338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2246_ _3476_/Q _2211_/B hold455/X _2201_/B _2214_/A vssd1 vssd1 vccd1 vccd1 _2246_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2177_ hold259/X _2587_/C _2176_/Y vssd1 vssd1 vccd1 vccd1 _2177_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_43_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput47 _2582_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_12
Xoutput58 _2473_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_12
XANTENNA__2878__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2912__S _2914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2030__A1 _2029_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2100_ _2108_/A _2100_/B vssd1 vssd1 vccd1 vccd1 _2100_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_27_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3080_ _3095_/A vssd1 vssd1 vccd1 vccd1 _3080_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2031_ hold832/X _2030_/X _2053_/S vssd1 vssd1 vccd1 vccd1 _2031_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2933_ _3055_/A vssd1 vssd1 vccd1 vccd1 _2933_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2864_ _2339_/B hold620/X _2864_/S vssd1 vssd1 vccd1 vccd1 _2864_/X sky130_fd_sc_hd__mux2_1
X_2795_ hold267/X _2805_/A1 _2803_/S vssd1 vssd1 vccd1 vccd1 _2795_/X sky130_fd_sc_hd__mux2_1
X_1815_ _1745_/B _1815_/B vssd1 vssd1 vccd1 vccd1 _1815_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_13_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1746_ _1813_/A _3555_/Q _1795_/B vssd1 vssd1 vccd1 vccd1 _1772_/B sky130_fd_sc_hd__or3b_4
Xhold302 _3220_/Q vssd1 vssd1 vccd1 vccd1 hold302/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold313 _3267_/Q vssd1 vssd1 vccd1 vccd1 hold313/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold324 _2669_/X vssd1 vssd1 vccd1 vccd1 _3202_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 _3256_/Q vssd1 vssd1 vccd1 vccd1 hold335/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 _3275_/Q vssd1 vssd1 vccd1 vccd1 hold368/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 _3444_/Q vssd1 vssd1 vccd1 vccd1 hold357/X sky130_fd_sc_hd__dlygate4sd3_1
X_1677_ hold65/X _1677_/B _1677_/C vssd1 vssd1 vccd1 vccd1 _2415_/A sky130_fd_sc_hd__and3_2
Xhold346 _2596_/X vssd1 vssd1 vccd1 vccd1 _3141_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 _2783_/X vssd1 vssd1 vccd1 vccd1 _3304_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3416_ _3416_/CLK _3416_/D vssd1 vssd1 vccd1 vccd1 _3416_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3347_ _3642_/CLK _3347_/D _2922_/Y vssd1 vssd1 vccd1 vccd1 _3347_/Q sky130_fd_sc_hd__dfrtp_1
Xhold1002 _2236_/X vssd1 vssd1 vccd1 vccd1 _3480_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1024 _2139_/X vssd1 vssd1 vccd1 vccd1 _3502_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 _2161_/X vssd1 vssd1 vccd1 vccd1 _3496_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1035 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 input13/A sky130_fd_sc_hd__dlygate4sd3_1
X_3278_ _3305_/CLK _3278_/D vssd1 vssd1 vccd1 vccd1 _3278_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1046 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 hold119/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1057 _3638_/Q vssd1 vssd1 vccd1 vccd1 hold207/A sky130_fd_sc_hd__dlygate4sd3_1
X_2229_ _2211_/B _2229_/B _2229_/C _2229_/D vssd1 vssd1 vccd1 vccd1 _2229_/X sky130_fd_sc_hd__and4b_1
XFILLER_0_63_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold880 _1800_/X vssd1 vssd1 vccd1 vccd1 _3559_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 _2328_/X vssd1 vssd1 vccd1 vccd1 hold891/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold937_A _3642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2907__S _2914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1600_ _2149_/A vssd1 vssd1 vccd1 vccd1 _1600_/Y sky130_fd_sc_hd__inv_2
X_2580_ _2580_/A hold29/A vssd1 vssd1 vccd1 vccd1 _2580_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1988__S1 _2044_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3201_ _3331_/CLK _3201_/D vssd1 vssd1 vccd1 vccd1 _3201_/Q sky130_fd_sc_hd__dfxtp_1
X_3132_ _3133_/A vssd1 vssd1 vccd1 vccd1 _3132_/Y sky130_fd_sc_hd__inv_2
X_3063_ _3065_/A vssd1 vssd1 vccd1 vccd1 _3063_/Y sky130_fd_sc_hd__inv_2
X_2014_ hold154/X hold185/X hold163/X hold148/X _1590_/A _2222_/A vssd1 vssd1 vccd1
+ vccd1 _2014_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2916_ _3437_/Q _1606_/Y _2915_/Y hold886/X vssd1 vssd1 vccd1 vccd1 _2916_/X sky130_fd_sc_hd__o2bb2a_1
X_2847_ _2101_/X hold686/X _2853_/S vssd1 vssd1 vccd1 vccd1 _2847_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold110 _2287_/X vssd1 vssd1 vccd1 vccd1 _2409_/B sky130_fd_sc_hd__dlygate4sd3_1
X_2778_ _2808_/A1 hold148/X _2783_/S vssd1 vssd1 vccd1 vccd1 _2778_/X sky130_fd_sc_hd__mux2_1
X_1729_ _3537_/Q _3454_/Q vssd1 vssd1 vccd1 vccd1 _1729_/Y sky130_fd_sc_hd__nand2b_1
Xhold121 _1674_/X vssd1 vssd1 vccd1 vccd1 _3608_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 _2677_/X vssd1 vssd1 vccd1 vccd1 _3209_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1979__S1 _2193_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold132 _3281_/Q vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 input20/X vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold165 _3297_/Q vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _3245_/Q vssd1 vssd1 vccd1 vccd1 hold154/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 _3306_/Q vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 _2407_/A vssd1 vssd1 vccd1 vccd1 _2419_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1631__S hold8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2637__S _2640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2701_ _2811_/A1 hold394/X _2703_/S vssd1 vssd1 vccd1 vccd1 _2701_/X sky130_fd_sc_hd__mux2_1
X_2632_ _2342_/B hold608/X _2640_/S vssd1 vssd1 vccd1 vccd1 _2632_/X sky130_fd_sc_hd__mux2_1
X_2563_ hold23/A hold7/A hold67/A _3593_/Q _2511_/Y vssd1 vssd1 vccd1 vccd1 _2563_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2401__A hold44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2494_ _3341_/Q _3588_/Q _2568_/C vssd1 vssd1 vccd1 vccd1 _2494_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2547__S _3522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3115_ _3121_/A vssd1 vssd1 vccd1 vccd1 _3115_/Y sky130_fd_sc_hd__inv_2
X_3046_ _3073_/A vssd1 vssd1 vccd1 vccd1 _3046_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2981__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout82 hold959/X vssd1 vssd1 vccd1 vccd1 _2905_/B sky130_fd_sc_hd__clkbuf_8
Xfanout71 _2096_/Y vssd1 vssd1 vccd1 vccd1 _2342_/B sky130_fd_sc_hd__buf_4
Xfanout93 _3489_/Q vssd1 vssd1 vccd1 vccd1 _2045_/S sky130_fd_sc_hd__buf_6
XFILLER_0_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2390__B1 _3341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3499_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1994_ _1985_/S _1994_/B vssd1 vssd1 vccd1 vccd1 _1994_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2615_ _2079_/A hold786/X _2618_/S vssd1 vssd1 vccd1 vccd1 _2615_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3595_ _3614_/CLK _3595_/D _3086_/Y vssd1 vssd1 vccd1 vccd1 _3595_/Q sky130_fd_sc_hd__dfrtp_1
X_2546_ _2545_/X _2544_/X _2551_/S vssd1 vssd1 vccd1 vccd1 _2546_/X sky130_fd_sc_hd__mux2_1
X_2477_ _3599_/Q _2568_/B _2417_/B _3343_/Q vssd1 vssd1 vccd1 vccd1 _2477_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3029_ _3036_/A vssd1 vssd1 vccd1 vccd1 _3029_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2531__S1 _1942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2047__S0 _1590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2675__A1 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold709 _2848_/X vssd1 vssd1 vccd1 vccd1 _3371_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2400_ hold52/X _2403_/B vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__and2_1
X_3380_ _3604_/CLK _3380_/D _2928_/Y vssd1 vssd1 vccd1 vccd1 _3380_/Q sky130_fd_sc_hd__dfrtp_1
X_2331_ _3381_/Q _2269_/X hold847/X vssd1 vssd1 vccd1 vccd1 _2331_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2262_ _2231_/D _2261_/X _1950_/B vssd1 vssd1 vccd1 vccd1 _2272_/C sky130_fd_sc_hd__a21oi_2
X_2193_ _2193_/A1 _2224_/B _2190_/A vssd1 vssd1 vccd1 vccd1 _2194_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout121_A _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1977_ _3513_/Q _1976_/Y _2052_/S vssd1 vssd1 vccd1 vccd1 _1977_/X sky130_fd_sc_hd__mux2_1
X_3578_ _3579_/CLK _3578_/D _3072_/Y vssd1 vssd1 vccd1 vccd1 _3578_/Q sky130_fd_sc_hd__dfrtp_1
X_2529_ _3185_/Q _3338_/Q _3167_/Q _3149_/Q _1911_/C _2550_/S1 vssd1 vssd1 vccd1 vccd1
+ _2529_/X sky130_fd_sc_hd__mux4_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__clkbuf_2
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 input8/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2820__A1 _2079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2880_ _2111_/B hold768/X _2884_/S vssd1 vssd1 vccd1 vccd1 _2880_/X sky130_fd_sc_hd__mux2_1
X_1900_ _3523_/Q _2598_/C vssd1 vssd1 vccd1 vccd1 _1902_/B sky130_fd_sc_hd__nand2_1
X_1831_ hold836/X _3545_/Q _1831_/S vssd1 vssd1 vccd1 vccd1 _1831_/X sky130_fd_sc_hd__mux2_1
X_1762_ hold977/X _2383_/C _1761_/X vssd1 vssd1 vccd1 vccd1 _1762_/X sky130_fd_sc_hd__o21a_1
X_1693_ _1707_/A _1707_/B vssd1 vssd1 vccd1 vccd1 _1705_/B sky130_fd_sc_hd__or2_1
Xhold517 _2872_/X vssd1 vssd1 vccd1 vccd1 _3398_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3501_ _3551_/CLK _3501_/D _2995_/Y vssd1 vssd1 vccd1 vccd1 _3501_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold506 _3591_/Q vssd1 vssd1 vccd1 vccd1 _2335_/A sky130_fd_sc_hd__dlygate4sd3_1
X_3432_ _3435_/CLK _3432_/D vssd1 vssd1 vccd1 vccd1 _3432_/Q sky130_fd_sc_hd__dfxtp_1
Xhold528 _3357_/Q vssd1 vssd1 vccd1 vccd1 hold528/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 _2868_/X vssd1 vssd1 vccd1 vccd1 _3394_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ _3414_/CLK _3363_/D vssd1 vssd1 vccd1 vccd1 _3363_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_41_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3427_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2431__S0 _1911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _3488_/CLK _3294_/D vssd1 vssd1 vccd1 vccd1 _3294_/Q sky130_fd_sc_hd__dfxtp_1
X_2314_ _2314_/A _2314_/B vssd1 vssd1 vccd1 vccd1 _2314_/Y sky130_fd_sc_hd__xnor2_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2245_ hold454/X _2242_/B _2243_/X _2244_/X vssd1 vssd1 vccd1 vccd1 _2245_/X sky130_fd_sc_hd__o211a_1
X_2176_ _2587_/C _2225_/B _2214_/A vssd1 vssd1 vccd1 vccd1 _2176_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2811__A1 _2811_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput48 _3650_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_12
Xoutput59 _3659_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_12
XANTENNA__1634__S hold8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2802__A1 _2812_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2869__A1 _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2030_ hold814/X _2029_/Y _2052_/S vssd1 vssd1 vccd1 vccd1 _2030_/X sky130_fd_sc_hd__mux2_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2932_ _3055_/A vssd1 vssd1 vccd1 vccd1 _2932_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2863_ _2338_/B hold794/X _2864_/S vssd1 vssd1 vccd1 vccd1 _2863_/X sky130_fd_sc_hd__mux2_1
X_1814_ _1813_/A _1810_/Y _1817_/B vssd1 vssd1 vccd1 vccd1 _1814_/X sky130_fd_sc_hd__a21o_1
X_2794_ _2794_/A _2794_/B _2794_/C vssd1 vssd1 vccd1 vccd1 _2803_/S sky130_fd_sc_hd__nor3_4
XFILLER_0_25_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1745_ _1813_/A _1745_/B _1795_/B vssd1 vssd1 vccd1 vccd1 _1745_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_0_80_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold325 _3265_/Q vssd1 vssd1 vccd1 vccd1 hold325/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 _2742_/X vssd1 vssd1 vccd1 vccd1 _3267_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold303 _2690_/X vssd1 vssd1 vccd1 vccd1 _3220_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 _3268_/Q vssd1 vssd1 vccd1 vccd1 hold347/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 _2751_/X vssd1 vssd1 vccd1 vccd1 _3275_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold358 _3201_/Q vssd1 vssd1 vccd1 vccd1 hold358/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 _2730_/X vssd1 vssd1 vccd1 vccd1 _3256_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2309__B1 _1996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1676_ hold18/X hold6/X vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__nor2_2
XFILLER_0_68_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3415_ _3416_/CLK _3415_/D vssd1 vssd1 vccd1 vccd1 _3415_/Q sky130_fd_sc_hd__dfxtp_1
X_3346_ _3580_/CLK _3346_/D _2921_/Y vssd1 vssd1 vccd1 vccd1 _3346_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1014 _3552_/Q vssd1 vssd1 vccd1 vccd1 _1580_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1003 hold1056/X vssd1 vssd1 vccd1 vccd1 _2149_/A sky130_fd_sc_hd__clkbuf_2
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1025 _3537_/Q vssd1 vssd1 vccd1 vccd1 _1849_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3277_ _3316_/CLK _3277_/D vssd1 vssd1 vccd1 vccd1 _3277_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1047 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 _3515_/Q vssd1 vssd1 vccd1 vccd1 hold499/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1036 _1625_/X vssd1 vssd1 vccd1 vccd1 _1626_/A sky130_fd_sc_hd__dlygate4sd3_1
X_2228_ _3490_/Q _2228_/B vssd1 vssd1 vccd1 vccd1 _2229_/D sky130_fd_sc_hd__or2_1
X_2159_ _2129_/A _2152_/Y _2158_/X vssd1 vssd1 vccd1 vccd1 _2159_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold870 _2330_/X vssd1 vssd1 vccd1 vccd1 _3382_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold881 _3500_/Q vssd1 vssd1 vccd1 vccd1 _2134_/C sky130_fd_sc_hd__clkbuf_2
Xhold892 _3574_/Q vssd1 vssd1 vccd1 vccd1 _1707_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2720__A0 _2810_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2787__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3200_ _3328_/CLK _3200_/D vssd1 vssd1 vccd1 vccd1 _3200_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2711__A0 _2811_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3131_ _3131_/A vssd1 vssd1 vccd1 vccd1 _3131_/Y sky130_fd_sc_hd__inv_2
X_3062_ _3065_/A vssd1 vssd1 vccd1 vccd1 _3062_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2013_ hold157/X _3281_/Q hold144/X hold150/X _1590_/A _2222_/A vssd1 vssd1 vccd1
+ vccd1 _2013_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2778__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2915_ _3055_/A _2915_/B _2915_/C vssd1 vssd1 vccd1 vccd1 _2915_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_5_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2846_ _2097_/A hold688/X _2853_/S vssd1 vssd1 vccd1 vccd1 _2846_/X sky130_fd_sc_hd__mux2_1
X_2777_ _2807_/A1 hold250/X _2783_/S vssd1 vssd1 vccd1 vccd1 _2777_/X sky130_fd_sc_hd__mux2_1
Xhold100 _3600_/Q vssd1 vssd1 vccd1 vccd1 hold100/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 input28/A sky130_fd_sc_hd__dlygate4sd3_1
X_1728_ _3540_/Q _3457_/Q vssd1 vssd1 vccd1 vccd1 _1728_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold111 _2441_/B vssd1 vssd1 vccd1 vccd1 _2585_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 _2758_/X vssd1 vssd1 vccd1 vccd1 _3281_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 _3272_/Q vssd1 vssd1 vccd1 vccd1 hold144/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 _2776_/X vssd1 vssd1 vccd1 vccd1 _3297_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 _2718_/X vssd1 vssd1 vccd1 vccd1 _3245_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1659_ _1659_/A hold26/X input9/X vssd1 vssd1 vccd1 vccd1 _1677_/B sky130_fd_sc_hd__and3_1
Xhold177 _2584_/X vssd1 vssd1 vccd1 vccd1 _3606_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _2786_/X vssd1 vssd1 vccd1 vccd1 _3306_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _1663_/X vssd1 vssd1 vccd1 vccd1 _1667_/S sky130_fd_sc_hd__clkbuf_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2702__A0 _2812_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _3331_/CLK _3329_/D vssd1 vssd1 vccd1 vccd1 _3329_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2769__A0 _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2979__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2700_ _2810_/A1 hold311/X _2703_/S vssd1 vssd1 vccd1 vccd1 _2700_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2631_ _3526_/Q _2905_/B _2875_/A vssd1 vssd1 vccd1 vccd1 _2640_/S sky130_fd_sc_hd__or3_4
X_2562_ _2506_/S _2552_/Y _2556_/X _2560_/X _2561_/Y vssd1 vssd1 vccd1 vccd1 _2562_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_10_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2493_ hold67/A _2568_/C vssd1 vssd1 vccd1 vccd1 _2493_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3114_ _3114_/A vssd1 vssd1 vccd1 vccd1 _3114_/Y sky130_fd_sc_hd__inv_2
X_3045_ _3121_/A vssd1 vssd1 vccd1 vccd1 _3045_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2829_ hold770/X _2111_/B _2833_/S vssd1 vssd1 vccd1 vccd1 _2829_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold196_A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1642__S hold8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout83 _1911_/A vssd1 vssd1 vccd1 vccd1 _2551_/S sky130_fd_sc_hd__buf_6
Xfanout72 _2091_/X vssd1 vssd1 vccd1 vccd1 _2097_/A sky130_fd_sc_hd__buf_4
XANTENNA__1965__A1 _1985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout94 _2193_/A1 vssd1 vssd1 vccd1 vccd1 _2044_/S1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2914__A0 _2339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_7_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1993_ _1992_/X _1991_/X _2045_/S vssd1 vssd1 vccd1 vccd1 _1994_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2614_ _2111_/B hold696/X _2618_/S vssd1 vssd1 vccd1 vccd1 _2614_/X sky130_fd_sc_hd__mux2_1
X_3594_ _3609_/CLK _3594_/D _3085_/Y vssd1 vssd1 vccd1 vccd1 _3594_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2545_ _3177_/Q _3426_/Q _3417_/Q _3159_/Q _2554_/S0 _1942_/A vssd1 vssd1 vccd1 vccd1
+ _2545_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_76_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2476_ _2476_/A _2476_/B vssd1 vssd1 vccd1 vccd1 _2476_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3028_ _3036_/A vssd1 vssd1 vccd1 vccd1 _3028_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2293__S hold30/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1947__A1 _3522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1637__S hold8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2047__S1 _2222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2468__S _2551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2330_ _1891_/A _3382_/Q hold869/X vssd1 vssd1 vccd1 vccd1 _2330_/X sky130_fd_sc_hd__o21ba_1
X_2261_ _2261_/A _2261_/B _2260_/X vssd1 vssd1 vccd1 vccd1 _2261_/X sky130_fd_sc_hd__or3b_1
X_2192_ _2189_/X _2242_/B _2191_/A _2196_/B vssd1 vssd1 vccd1 vccd1 _2192_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1976_ _1976_/A vssd1 vssd1 vccd1 vccd1 _1976_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3577_ _3579_/CLK _3577_/D _3071_/Y vssd1 vssd1 vccd1 vccd1 _3577_/Q sky130_fd_sc_hd__dfrtp_1
X_2528_ _3407_/Q _3398_/Q _3389_/Q _3434_/Q _1911_/C _2550_/S1 vssd1 vssd1 vccd1 vccd1
+ _2528_/X sky130_fd_sc_hd__mux4_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ _3609_/Q _2441_/A _2458_/X vssd1 vssd1 vccd1 vccd1 _2459_/X sky130_fd_sc_hd__a21o_1
Xhold26 input8/X vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2751__S _2753_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2593__A1 _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1830_ hold859/X hold836/X _1831_/S vssd1 vssd1 vccd1 vccd1 _1830_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2027__A_N _1985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3500_ _3551_/CLK _3500_/D _2994_/Y vssd1 vssd1 vccd1 vccd1 _3500_/Q sky130_fd_sc_hd__dfrtp_1
X_1761_ _1811_/A _1761_/B _1772_/B vssd1 vssd1 vccd1 vccd1 _1761_/X sky130_fd_sc_hd__or3_1
X_1692_ _1692_/A _1692_/B _1711_/B vssd1 vssd1 vccd1 vccd1 _1707_/B sky130_fd_sc_hd__or3_1
Xhold518 _3400_/Q vssd1 vssd1 vccd1 vccd1 hold518/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold507 _2335_/Y vssd1 vssd1 vccd1 vccd1 _3379_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold529 _2832_/X vssd1 vssd1 vccd1 vccd1 _3357_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3431_ _3433_/CLK _3431_/D vssd1 vssd1 vccd1 vccd1 _3431_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ _3423_/CLK _3362_/D vssd1 vssd1 vccd1 vccd1 _3362_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2431__S1 _1942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2313_ _1565_/Y _1976_/A _1985_/X _2312_/Y vssd1 vssd1 vccd1 vccd1 _2314_/B sky130_fd_sc_hd__o31a_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _3610_/CLK _3293_/D vssd1 vssd1 vccd1 vccd1 _3293_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ _2794_/B _2244_/B vssd1 vssd1 vccd1 vccd1 _2244_/X sky130_fd_sc_hd__xor2_1
X_2175_ _2175_/A _2175_/B vssd1 vssd1 vccd1 vccd1 _2225_/B sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3318_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1959_ hold457/X hold450/X hold404/X hold418/X _2044_/S0 _2044_/S1 vssd1 vssd1 vccd1
+ vccd1 _1959_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_31_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3629_ _3629_/CLK hold81/X _3120_/Y vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__dfrtp_1
Xoutput38 _2391_/X vssd1 vssd1 vccd1 vccd1 uart_irq sky130_fd_sc_hd__buf_12
Xoutput49 _3651_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_12
XANTENNA__2746__S _2753_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2931_ _3055_/A vssd1 vssd1 vccd1 vccd1 _2931_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_84_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2862_ _2075_/B hold578/X _2864_/S vssd1 vssd1 vccd1 vccd1 _2862_/X sky130_fd_sc_hd__mux2_1
X_2793_ _2813_/A1 hold349/X _2793_/S vssd1 vssd1 vccd1 vccd1 _2793_/X sky130_fd_sc_hd__mux2_1
X_1813_ _1813_/A _1817_/B vssd1 vssd1 vccd1 vccd1 _1813_/Y sky130_fd_sc_hd__nor2_1
X_1744_ _1744_/A _3553_/Q _3552_/Q vssd1 vssd1 vccd1 vccd1 _1813_/A sky130_fd_sc_hd__nand3_2
Xhold326 _2740_/X vssd1 vssd1 vccd1 vccd1 _3265_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold304 _3598_/Q vssd1 vssd1 vccd1 vccd1 hold304/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold52_A hold52/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold315 _3238_/Q vssd1 vssd1 vccd1 vccd1 hold315/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 _2743_/X vssd1 vssd1 vccd1 vccd1 _3268_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1675_ _2585_/A _3607_/Q _1675_/S vssd1 vssd1 vccd1 vccd1 _1675_/X sky130_fd_sc_hd__mux2_1
Xhold337 _3310_/Q vssd1 vssd1 vccd1 vccd1 hold337/X sky130_fd_sc_hd__dlygate4sd3_1
X_3414_ _3414_/CLK _3414_/D vssd1 vssd1 vccd1 vccd1 _3414_/Q sky130_fd_sc_hd__dfxtp_1
Xhold359 _2668_/X vssd1 vssd1 vccd1 vccd1 _3201_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3345_ _3580_/CLK _3345_/D _2920_/Y vssd1 vssd1 vccd1 vccd1 _3345_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3276_ _3316_/CLK _3276_/D vssd1 vssd1 vccd1 vccd1 _3276_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1015 _1820_/Y vssd1 vssd1 vccd1 vccd1 _1821_/B1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1004 _2368_/Y vssd1 vssd1 vccd1 vccd1 _3346_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1037 _3578_/Q vssd1 vssd1 vccd1 vccd1 _1697_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 _3558_/Q vssd1 vssd1 vccd1 vccd1 _1797_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ _3490_/Q _2228_/B vssd1 vssd1 vccd1 vccd1 _2229_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_84_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1059 _3572_/Q vssd1 vssd1 vccd1 vccd1 hold818/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2158_ _1951_/Y _2130_/C _2149_/X _2161_/S vssd1 vssd1 vccd1 vccd1 _2158_/X sky130_fd_sc_hd__a31o_1
X_2089_ _3546_/Q _2089_/B vssd1 vssd1 vccd1 vccd1 _2089_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__2796__A1 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2548__B2 _2506_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2548__A1 _2583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold860 _1830_/X vssd1 vssd1 vccd1 vccd1 _3546_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 _3439_/Q vssd1 vssd1 vccd1 vccd1 _1824_/A sky130_fd_sc_hd__buf_2
Xhold882 _2144_/Y vssd1 vssd1 vccd1 vccd1 _3500_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout94_A _2193_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold893 _1707_/Y vssd1 vssd1 vccd1 vccd1 hold893/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2224__B _2224_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3130_ _3133_/A vssd1 vssd1 vccd1 vccd1 _3130_/Y sky130_fd_sc_hd__inv_2
X_3061_ _3065_/A vssd1 vssd1 vccd1 vccd1 _3061_/Y sky130_fd_sc_hd__inv_2
X_2012_ _2010_/X _2011_/X _2045_/S vssd1 vssd1 vccd1 vccd1 _2012_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2914_ _2339_/B hold618/X _2914_/S vssd1 vssd1 vccd1 vccd1 _2914_/X sky130_fd_sc_hd__mux2_1
X_2845_ _2342_/B hold660/X _2853_/S vssd1 vssd1 vccd1 vccd1 _2845_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2776_ _2806_/A1 hold165/X _2783_/S vssd1 vssd1 vccd1 vccd1 _2776_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold101 _3450_/Q vssd1 vssd1 vccd1 vccd1 _1720_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 input28/X vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_79_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1727_ _1582_/Y _3459_/Q _3453_/Q _1847_/A vssd1 vssd1 vccd1 vccd1 _1735_/A sky130_fd_sc_hd__o22ai_1
XFILLER_0_13_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold134 _3236_/Q vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 _2585_/X vssd1 vssd1 vccd1 vccd1 _3595_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _2748_/X vssd1 vssd1 vccd1 vccd1 _3272_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 _3288_/Q vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 wbs_we_i vssd1 vssd1 vccd1 vccd1 input37/A sky130_fd_sc_hd__dlygate4sd3_1
X_1658_ hold18/X _1658_/B vssd1 vssd1 vccd1 vccd1 _2410_/A sky130_fd_sc_hd__nor2_2
Xhold189 _3279_/Q vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 _3261_/Q vssd1 vssd1 vccd1 vccd1 hold178/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3328_ _3328_/CLK _3328_/D vssd1 vssd1 vccd1 vccd1 _3328_/Q sky130_fd_sc_hd__dfxtp_1
X_1589_ _1589_/A vssd1 vssd1 vccd1 vccd1 _2130_/A sky130_fd_sc_hd__inv_2
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ _3513_/CLK _3259_/D vssd1 vssd1 vccd1 vccd1 _3259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold690 _3179_/Q vssd1 vssd1 vccd1 vccd1 hold690/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2630_ _3524_/Q _3523_/Q _2630_/C vssd1 vssd1 vccd1 vccd1 _2875_/A sky130_fd_sc_hd__or3_2
XFILLER_0_54_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2561_ _1595_/Y _2511_/B _2506_/S vssd1 vssd1 vccd1 vccd1 _2561_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2492_ _3341_/Q _1678_/X _2412_/Y _3600_/Q vssd1 vssd1 vccd1 vccd1 _2492_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_10_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2696__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3113_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3113_/Y sky130_fd_sc_hd__inv_2
X_3044_ _3044_/A vssd1 vssd1 vccd1 vccd1 _3044_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_81_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2828_ hold548/X _2105_/B _2833_/S vssd1 vssd1 vccd1 vccd1 _2828_/X sky130_fd_sc_hd__mux2_1
X_2759_ hold384/X _2809_/A1 _2763_/S vssd1 vssd1 vccd1 vccd1 _2759_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2687__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2611__A0 _2097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout73 _2081_/X vssd1 vssd1 vccd1 vccd1 _2339_/B sky130_fd_sc_hd__buf_4
Xfanout95 _2193_/A1 vssd1 vssd1 vccd1 vccd1 _2222_/A sky130_fd_sc_hd__clkbuf_8
Xfanout84 _1942_/A vssd1 vssd1 vccd1 vccd1 _2550_/S1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2664__S _2672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1653__A1 _2397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1992_ _3247_/Q _3319_/Q _3310_/Q _3301_/Q _1590_/A _2222_/A vssd1 vssd1 vccd1 vccd1
+ _1992_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2602__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_35_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3576_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3593_ _3633_/CLK hold15/X _3084_/Y vssd1 vssd1 vccd1 vccd1 _3593_/Q sky130_fd_sc_hd__dfrtp_1
X_2613_ _2105_/B hold802/X _2618_/S vssd1 vssd1 vccd1 vccd1 _2613_/X sky130_fd_sc_hd__mux2_1
X_2544_ _3375_/Q _3357_/Q _3366_/Q _3195_/Q _2554_/S0 _1911_/B vssd1 vssd1 vccd1 vccd1
+ _2544_/X sky130_fd_sc_hd__mux4_1
X_2475_ _3614_/Q _2439_/A _2406_/X vssd1 vssd1 vccd1 vccd1 _2475_/X sky130_fd_sc_hd__a21o_1
XANTENNA__2669__A0 _2810_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2516__S0 _1943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3027_ _3036_/A vssd1 vssd1 vccd1 vccd1 _3027_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2841__A0 _2075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1644__A1 _2585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2749__S _2753_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1889__A _2231_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1635__A1 hold14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2260_ _2260_/A _2260_/B _3477_/Q vssd1 vssd1 vccd1 vccd1 _2260_/X sky130_fd_sc_hd__and3_1
X_2191_ _2191_/A _2194_/A vssd1 vssd1 vccd1 vccd1 _2242_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1975_ _1985_/S _1970_/X _1974_/X vssd1 vssd1 vccd1 vccd1 _1976_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_28_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3576_ _3576_/CLK _3576_/D _3070_/Y vssd1 vssd1 vccd1 vccd1 _3576_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout107_A hold126/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2527_ _2511_/Y _2525_/X _2526_/X _2511_/B _3450_/Q vssd1 vssd1 vccd1 vccd1 _2527_/X
+ sky130_fd_sc_hd__a32o_1
X_2458_ _3586_/Q hold67/A _2508_/B _2457_/X vssd1 vssd1 vccd1 vccd1 _2458_/X sky130_fd_sc_hd__o211a_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ _3596_/Q _3594_/Q _3342_/Q _3598_/Q _2386_/X vssd1 vssd1 vccd1 vccd1 _2391_/B
+ sky130_fd_sc_hd__a221o_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1891__B _2231_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1760_ hold975/X _2383_/C _1759_/X vssd1 vssd1 vccd1 vccd1 _1760_/X sky130_fd_sc_hd__o21a_1
X_1691_ _3594_/Q _3476_/Q hold857/X vssd1 vssd1 vccd1 vccd1 _1691_/X sky130_fd_sc_hd__o21ba_1
Xhold508 _3590_/Q vssd1 vssd1 vccd1 vccd1 _2337_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3430_ _3435_/CLK _3430_/D vssd1 vssd1 vccd1 vccd1 _3430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold519 _2874_/X vssd1 vssd1 vccd1 vccd1 _3400_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2336__A2 _1889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3361_ _3369_/CLK _3361_/D vssd1 vssd1 vccd1 vccd1 _3361_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2312_ _1565_/Y _1976_/A _1985_/X _2311_/X vssd1 vssd1 vccd1 vccd1 _2312_/Y sky130_fd_sc_hd__o211ai_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ _3305_/CLK _3292_/D vssd1 vssd1 vccd1 vccd1 _3292_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2243_ _2226_/A _2243_/B _2243_/C _2243_/D vssd1 vssd1 vccd1 vccd1 _2243_/X sky130_fd_sc_hd__and4b_1
XFILLER_0_73_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2174_ _3492_/Q _3491_/Q _2794_/B vssd1 vssd1 vccd1 vccd1 _2175_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1958_ hold442/X hold452/X hold436/X hold440/X _2044_/S0 _2044_/S1 vssd1 vssd1 vccd1
+ vccd1 _1958_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1889_ _2231_/D vssd1 vssd1 vccd1 vccd1 _1889_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3628_ _3629_/CLK _3628_/D _3119_/Y vssd1 vssd1 vccd1 vccd1 _3628_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput39 _3443_/Q vssd1 vssd1 vccd1 vccd1 uart_tx sky130_fd_sc_hd__buf_12
XANTENNA__2327__A2 _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3559_ _3559_/CLK _3559_/D _3053_/Y vssd1 vssd1 vccd1 vccd1 _3559_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2762__S _2763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2930_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2930_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2672__S _2672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2861_ _2079_/A hold718/X _2864_/S vssd1 vssd1 vccd1 vccd1 _2861_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2006__A1 _1985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2792_ _2812_/A1 hold276/X _2793_/S vssd1 vssd1 vccd1 vccd1 _2792_/X sky130_fd_sc_hd__mux2_1
X_1812_ _1811_/A _1810_/Y _1811_/Y _1795_/B vssd1 vssd1 vccd1 vccd1 _1817_/B sky130_fd_sc_hd__o211ai_4
XFILLER_0_4_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1743_ _1743_/A _1743_/B _1743_/C wire80/X vssd1 vssd1 vccd1 vccd1 _2381_/A sky130_fd_sc_hd__nor4b_4
Xhold305 _3247_/Q vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
X_1674_ _2395_/A _3608_/Q _1675_/S vssd1 vssd1 vccd1 vccd1 _1674_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold316 _2710_/X vssd1 vssd1 vccd1 vccd1 _3238_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 _3313_/Q vssd1 vssd1 vccd1 vccd1 hold349/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 _2790_/X vssd1 vssd1 vccd1 vccd1 _3310_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3413_ _3423_/CLK _3413_/D vssd1 vssd1 vccd1 vccd1 _3413_/Q sky130_fd_sc_hd__dfxtp_1
Xhold327 _3204_/Q vssd1 vssd1 vccd1 vccd1 hold327/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3344_ _3642_/CLK _3344_/D _2919_/Y vssd1 vssd1 vccd1 vccd1 _3344_/Q sky130_fd_sc_hd__dfstp_1
X_3275_ _3319_/CLK _3275_/D vssd1 vssd1 vccd1 vccd1 _3275_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1005 _3553_/Q vssd1 vssd1 vccd1 vccd1 _1774_/C sky130_fd_sc_hd__dlygate4sd3_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1038 _3464_/Q vssd1 vssd1 vccd1 vccd1 _2263_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1027 _3465_/Q vssd1 vssd1 vccd1 vccd1 _1592_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 _1821_/X vssd1 vssd1 vccd1 vccd1 _3553_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ _2226_/A _2243_/B _2243_/C _2226_/D vssd1 vssd1 vccd1 vccd1 _2229_/B sky130_fd_sc_hd__and4_1
XFILLER_0_84_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2157_ _2161_/S _2156_/Y hold952/X vssd1 vssd1 vccd1 vccd1 _2157_/X sky130_fd_sc_hd__o21a_1
X_2088_ _2121_/A _2088_/B vssd1 vssd1 vccd1 vccd1 _2088_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_63_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1661__A_N hold65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold850 _2239_/X vssd1 vssd1 vccd1 vccd1 _3478_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 _3548_/Q vssd1 vssd1 vccd1 vccd1 hold861/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 _1831_/S vssd1 vssd1 vccd1 vccd1 _1833_/S sky130_fd_sc_hd__clkbuf_2
Xhold894 _1708_/Y vssd1 vssd1 vccd1 vccd1 _3574_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout87_A _1911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold883 hold883/A vssd1 vssd1 vccd1 vccd1 _2145_/D sky130_fd_sc_hd__buf_1
XANTENNA__2757__S _2763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2667__S _2672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3060_ _3065_/A vssd1 vssd1 vccd1 vccd1 _3060_/Y sky130_fd_sc_hd__inv_2
X_2011_ hold130/X hold142/X hold146/X hold140/X _2044_/S0 _2044_/S1 vssd1 vssd1 vccd1
+ vccd1 _2011_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2913_ _2338_/B hold798/X _2914_/S vssd1 vssd1 vccd1 vccd1 _2913_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2844_ _2875_/A _3526_/Q _2905_/B vssd1 vssd1 vccd1 vccd1 _2853_/S sky130_fd_sc_hd__or3b_4
X_2775_ _2805_/A1 hold221/X _2783_/S vssd1 vssd1 vccd1 vccd1 _2775_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold124 _1673_/X vssd1 vssd1 vccd1 vccd1 _3609_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1726_ hold46/A _3538_/Q vssd1 vssd1 vccd1 vccd1 _1726_/X sky130_fd_sc_hd__and2b_1
Xhold113 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 input10/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _2708_/X vssd1 vssd1 vccd1 vccd1 _3236_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 _2301_/X vssd1 vssd1 vccd1 vccd1 _3450_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _2766_/X vssd1 vssd1 vccd1 vccd1 _3288_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 _3200_/Q vssd1 vssd1 vccd1 vccd1 hold146/X sky130_fd_sc_hd__dlygate4sd3_1
X_1657_ _1657_/A hold57/X _1657_/C hold5/X vssd1 vssd1 vccd1 vccd1 _1658_/B sky130_fd_sc_hd__or4b_2
Xhold157 _3290_/Q vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 _2736_/X vssd1 vssd1 vccd1 vccd1 _3261_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1588_ _1588_/A vssd1 vssd1 vccd1 vccd1 _1588_/Y sky130_fd_sc_hd__inv_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3327_ _3331_/CLK _3327_/D vssd1 vssd1 vccd1 vccd1 _3327_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _3493_/CLK _3258_/D vssd1 vssd1 vccd1 vccd1 _3258_/Q sky130_fd_sc_hd__dfxtp_1
X_2209_ _2212_/C _2209_/B vssd1 vssd1 vccd1 vccd1 _2216_/B sky130_fd_sc_hd__and2_1
X_3189_ _3369_/CLK _3189_/D vssd1 vssd1 vccd1 vccd1 _3189_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2010__S0 _2044_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold680 _3396_/Q vssd1 vssd1 vccd1 vccd1 hold680/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold691 _2642_/X vssd1 vssd1 vccd1 vccd1 _3179_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2560_ hold54/A _2571_/B _2511_/B _2559_/X vssd1 vssd1 vccd1 vccd1 _2560_/X sky130_fd_sc_hd__a211o_1
X_2491_ _2506_/S _2490_/X _2483_/X vssd1 vssd1 vccd1 vccd1 _2491_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3112_ _3114_/A vssd1 vssd1 vccd1 vccd1 _3112_/Y sky130_fd_sc_hd__inv_2
X_3043_ _3073_/A vssd1 vssd1 vccd1 vccd1 _3043_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2860__S _2864_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2827_ hold532/X _2105_/A _2833_/S vssd1 vssd1 vccd1 vccd1 _2827_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2758_ hold132/X _2808_/A1 _2763_/S vssd1 vssd1 vccd1 vccd1 _2758_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1709_ _1692_/A _1711_/B _1692_/B vssd1 vssd1 vccd1 vccd1 _1709_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2689_ _2809_/A1 hold362/X _2693_/S vssd1 vssd1 vccd1 vccd1 _2689_/X sky130_fd_sc_hd__mux2_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_5_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3513_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2770__S _2773_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout74 _2076_/X vssd1 vssd1 vccd1 vccd1 _2338_/B sky130_fd_sc_hd__buf_4
Xfanout96 _3488_/Q vssd1 vssd1 vccd1 vccd1 _2193_/A1 sky130_fd_sc_hd__buf_4
Xfanout85 _1942_/A vssd1 vssd1 vccd1 vccd1 _1911_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__2470__S0 _2554_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2678__A1 _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1991_ _3292_/Q _3283_/Q _3274_/Q _3265_/Q _1590_/A _2222_/A vssd1 vssd1 vccd1 vccd1
+ _1991_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2680__S _2682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3077__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2612_ _2105_/A hold760/X _2618_/S vssd1 vssd1 vccd1 vccd1 _2612_/X sky130_fd_sc_hd__mux2_1
X_3592_ _3604_/CLK _3592_/D _3083_/Y vssd1 vssd1 vccd1 vccd1 _3592_/Q sky130_fd_sc_hd__dfrtp_1
X_2543_ _2542_/X _2541_/X _2551_/S vssd1 vssd1 vccd1 vccd1 _2543_/X sky130_fd_sc_hd__mux2_1
X_2474_ _3618_/Q _1645_/Y _2571_/B vssd1 vssd1 vccd1 vccd1 _2474_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_78_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3026_ _3036_/A vssd1 vssd1 vccd1 vccd1 _3026_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2516__S1 _2550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2452__S0 _2554_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2765__S _2773_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2832__A1 _2338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2899__A1 _2104_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2190_ _2190_/A _2222_/A _2224_/B vssd1 vssd1 vccd1 vccd1 _2194_/A sky130_fd_sc_hd__and3_1
XANTENNA__2675__S _2682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2823__A1 _2339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1974_ _2191_/A _1974_/B vssd1 vssd1 vccd1 vccd1 _1974_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3575_ _3576_/CLK _3575_/D _3069_/Y vssd1 vssd1 vccd1 vccd1 _3575_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2526_ hold87/A _1645_/Y _2568_/D _2524_/X vssd1 vssd1 vccd1 vccd1 _2526_/X sky130_fd_sc_hd__a22o_1
X_2457_ _3598_/Q _2568_/B _2417_/B _3342_/Q vssd1 vssd1 vccd1 vccd1 _2457_/X sky130_fd_sc_hd__o22a_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__buf_2
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
X_2388_ _3605_/Q _3381_/Q _3378_/Q hold78/A vssd1 vssd1 vccd1 vccd1 _2388_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3009_ _3114_/A vssd1 vssd1 vccd1 vccd1 _3009_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2750__A0 _2810_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2805__A1 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1690_ hold254/X _2585_/A hold21/X vssd1 vssd1 vccd1 vccd1 _3596_/D sky130_fd_sc_hd__mux2_1
Xhold509 _2337_/Y vssd1 vssd1 vccd1 vccd1 _3378_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3360_ _3369_/CLK _3360_/D vssd1 vssd1 vccd1 vccd1 _3360_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2741__A0 _2811_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2311_ _3626_/Q _3625_/Q _3624_/Q _3627_/Q vssd1 vssd1 vccd1 vccd1 _2311_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_57_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _3330_/CLK _3291_/D vssd1 vssd1 vccd1 vccd1 _3291_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2242_ _2794_/A _2242_/B vssd1 vssd1 vccd1 vccd1 _2243_/D sky130_fd_sc_hd__nand2_1
X_2173_ _2661_/B _2228_/B _2172_/Y _2214_/A vssd1 vssd1 vccd1 vccd1 _2173_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_0_25_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1957_ _3346_/Q _3344_/Q _1955_/Y _2375_/A vssd1 vssd1 vccd1 vccd1 _2053_/S sky130_fd_sc_hd__o211a_4
X_1888_ _2381_/A _1888_/B vssd1 vssd1 vccd1 vccd1 _2231_/D sky130_fd_sc_hd__nand2_4
XFILLER_0_24_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3627_ _3631_/CLK _3627_/D _3118_/Y vssd1 vssd1 vccd1 vccd1 _3627_/Q sky130_fd_sc_hd__dfstp_2
X_3558_ _3559_/CLK _3558_/D _3052_/Y vssd1 vssd1 vccd1 vccd1 _3558_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2732__A0 _2812_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2509_ _3589_/Q hold67/A vssd1 vssd1 vccd1 vccd1 _2509_/X sky130_fd_sc_hd__or2_1
X_3489_ _3610_/CLK _3489_/D _2983_/Y vssd1 vssd1 vccd1 vccd1 _3489_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_66_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2723__A0 _2813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2860_ _2111_/B hold714/X _2864_/S vssd1 vssd1 vccd1 vccd1 _2860_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1811_ _1811_/A _2111_/A vssd1 vssd1 vccd1 vccd1 _1811_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2791_ _2811_/A1 hold372/X _2793_/S vssd1 vssd1 vccd1 vccd1 _2791_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1742_ _2231_/B wire80/X vssd1 vssd1 vccd1 vccd1 _1950_/B sky130_fd_sc_hd__nand2_2
X_1673_ _2396_/A _3609_/Q _1675_/S vssd1 vssd1 vccd1 vccd1 _1673_/X sky130_fd_sc_hd__mux2_1
Xhold306 _2720_/X vssd1 vssd1 vccd1 vccd1 _3247_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 _3302_/Q vssd1 vssd1 vccd1 vccd1 hold317/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3412_ _3582_/CLK _3412_/D vssd1 vssd1 vccd1 vccd1 _3412_/Q sky130_fd_sc_hd__dfxtp_1
Xhold328 _2671_/X vssd1 vssd1 vccd1 vccd1 _3204_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 _3273_/Q vssd1 vssd1 vccd1 vccd1 hold339/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _3614_/CLK _3343_/D _2918_/Y vssd1 vssd1 vccd1 vccd1 _3343_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _3305_/CLK _3274_/D vssd1 vssd1 vccd1 vccd1 _3274_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1006 _1775_/B vssd1 vssd1 vccd1 vccd1 _1794_/A3 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1028 _2275_/Y vssd1 vssd1 vccd1 vccd1 _2276_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 _3474_/Q vssd1 vssd1 vccd1 vccd1 _2252_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 _3557_/Q vssd1 vssd1 vccd1 vccd1 _1797_/B sky130_fd_sc_hd__buf_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ _3489_/Q _2225_/B vssd1 vssd1 vccd1 vccd1 _2226_/D sky130_fd_sc_hd__xor2_1
X_2156_ _2156_/A _2156_/B vssd1 vssd1 vccd1 vccd1 _2156_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2863__S _2864_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2087_ _3547_/Q _2089_/B vssd1 vssd1 vccd1 vccd1 _2088_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2989_ _3120_/A vssd1 vssd1 vccd1 vccd1 _2989_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_31_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold840 _3479_/Q vssd1 vssd1 vccd1 vccd1 _2260_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 _3578_/Q vssd1 vssd1 vccd1 vccd1 _1700_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 _1829_/X vssd1 vssd1 vccd1 vccd1 _3547_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 _1825_/X vssd1 vssd1 vccd1 vccd1 _3551_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2705__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold895 _3461_/Q vssd1 vssd1 vccd1 vccd1 _2272_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold884 _2377_/X vssd1 vssd1 vccd1 vccd1 _3349_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2773__S _2773_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1995__A1 _1985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2010_ hold128/X hold136/X hold134/X hold138/X _2044_/S0 _2044_/S1 vssd1 vssd1 vccd1
+ vccd1 _2010_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_29_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3642_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2912_ _2075_/B hold604/X _2914_/S vssd1 vssd1 vccd1 vccd1 _2912_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2843_ _2339_/B hold736/X _2843_/S vssd1 vssd1 vccd1 vccd1 _2843_/X sky130_fd_sc_hd__mux2_1
X_2774_ _2794_/A _2794_/B _2804_/A vssd1 vssd1 vccd1 vccd1 _2783_/S sky130_fd_sc_hd__or3_4
XFILLER_0_79_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1725_ _3532_/Q hold72/X vssd1 vssd1 vccd1 vccd1 _1725_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_53_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold103 _3636_/Q vssd1 vssd1 vccd1 vccd1 _2263_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 input29/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 _2287_/A vssd1 vssd1 vccd1 vccd1 _1657_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 _2768_/X vssd1 vssd1 vccd1 vccd1 _3290_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _2667_/X vssd1 vssd1 vccd1 vccd1 _3200_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 _3137_/Q vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlygate4sd3_1
X_1656_ _2342_/A _2585_/A hold60/X vssd1 vssd1 vccd1 vccd1 _3615_/D sky130_fd_sc_hd__mux2_1
XANTENNA__2858__S _2864_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1587_ _1893_/A vssd1 vssd1 vccd1 vccd1 _2824_/B sky130_fd_sc_hd__inv_2
Xhold169 _3207_/Q vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _3328_/CLK _3326_/D vssd1 vssd1 vccd1 vccd1 _3326_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _3612_/CLK _3257_/D vssd1 vssd1 vccd1 vccd1 _3257_/Q sky130_fd_sc_hd__dfxtp_1
X_2208_ _2208_/A _2211_/B vssd1 vssd1 vccd1 vccd1 _2209_/B sky130_fd_sc_hd__or2_1
X_3188_ _3403_/CLK _3188_/D vssd1 vssd1 vccd1 vccd1 _3188_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2010__S1 _2044_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1674__A0 _2395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2139_ _2139_/A _2139_/B vssd1 vssd1 vccd1 vccd1 _2139_/X sky130_fd_sc_hd__and2_1
XFILLER_0_76_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold496_A _2200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold681 _2870_/X vssd1 vssd1 vccd1 vccd1 _3396_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold670 _3410_/Q vssd1 vssd1 vccd1 vccd1 hold670/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2768__S _2773_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold692 _3182_/Q vssd1 vssd1 vccd1 vccd1 hold692/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2008__S _2052_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2490_ _2489_/X _2486_/X _3522_/Q vssd1 vssd1 vccd1 vccd1 _2490_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2678__S _2682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3111_ _3114_/A vssd1 vssd1 vccd1 vccd1 _3111_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_65_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3042_ _3073_/A vssd1 vssd1 vccd1 vccd1 _3042_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1611__A _1660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2145__C _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2826_ hold526/X _2097_/A _2833_/S vssd1 vssd1 vccd1 vccd1 _2826_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2908__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2757_ hold280/X _2807_/A1 _2763_/S vssd1 vssd1 vccd1 vccd1 _2757_/X sky130_fd_sc_hd__mux2_1
X_1708_ _1705_/B hold893/X _3466_/D vssd1 vssd1 vccd1 vccd1 _1708_/Y sky130_fd_sc_hd__a21oi_1
X_2688_ _2808_/A1 hold130/X _2693_/S vssd1 vssd1 vccd1 vccd1 _2688_/X sky130_fd_sc_hd__mux2_1
X_1639_ hold80/X hold33/X hold8/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__mux2_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ _3493_/CLK _3309_/D vssd1 vssd1 vccd1 vccd1 _3309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout86 _3520_/Q vssd1 vssd1 vccd1 vccd1 _1942_/A sky130_fd_sc_hd__buf_4
Xfanout75 _2074_/X vssd1 vssd1 vccd1 vccd1 _2075_/B sky130_fd_sc_hd__buf_4
Xfanout97 _2224_/B vssd1 vssd1 vccd1 vccd1 _2044_/S0 sky130_fd_sc_hd__buf_8
XFILLER_0_64_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2470__S1 _1911_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1990_ _1988_/X _1989_/X _2045_/S vssd1 vssd1 vccd1 vccd1 _1990_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2611_ _2097_/A hold568/X _2618_/S vssd1 vssd1 vccd1 vccd1 _2611_/X sky130_fd_sc_hd__mux2_1
X_3591_ _3604_/CLK hold45/X _3082_/Y vssd1 vssd1 vccd1 vccd1 _3591_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2542_ _3186_/Q _3339_/Q _3168_/Q _3150_/Q _1943_/B _2550_/S1 vssd1 vssd1 vccd1 vccd1
+ _2542_/X sky130_fd_sc_hd__mux4_1
X_2473_ _2506_/S _2472_/X _2465_/X vssd1 vssd1 vccd1 vccd1 _2473_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_44_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3403_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1972__S0 _1590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3025_ _3036_/A vssd1 vssd1 vccd1 vccd1 _3025_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2809_ hold398/X _2809_/A1 _2813_/S vssd1 vssd1 vccd1 vccd1 _2809_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2452__S1 _1911_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2596__A1 _2812_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output43_A _2573_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2691__S _2693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1973_ _1972_/X _1971_/X _2045_/S vssd1 vssd1 vccd1 vccd1 _1974_/B sky130_fd_sc_hd__mux2_1
X_3574_ _3576_/CLK _3574_/D _3068_/Y vssd1 vssd1 vccd1 vccd1 _3574_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2525_ hold90/A hold7/A vssd1 vssd1 vccd1 vccd1 _2525_/X sky130_fd_sc_hd__or2_1
X_2456_ _3640_/Q _2511_/A _2511_/B vssd1 vssd1 vccd1 vccd1 _2456_/X sky130_fd_sc_hd__a21o_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 hold94/X vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2387_ hold68/A _3379_/Q _3343_/Q _3599_/Q vssd1 vssd1 vccd1 vccd1 _2391_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_78_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3008_ _3114_/A vssd1 vssd1 vccd1 vccd1 _3008_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_66_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2077__A _2338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2310_ _2310_/A _2310_/B vssd1 vssd1 vccd1 vccd1 _2314_/A sky130_fd_sc_hd__xnor2_1
X_3290_ _3318_/CLK _3290_/D vssd1 vssd1 vccd1 vccd1 _3290_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2686__S _2693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2241_ _2241_/A _2241_/B vssd1 vssd1 vccd1 vccd1 _2241_/Y sky130_fd_sc_hd__nor2_1
X_2172_ _2794_/A _2661_/B vssd1 vssd1 vccd1 vccd1 _2172_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1956_ _1956_/A _1956_/B vssd1 vssd1 vccd1 vccd1 _2375_/A sky130_fd_sc_hd__nand2_1
X_1887_ _2383_/A _1602_/Y _2915_/B vssd1 vssd1 vccd1 vccd1 _1888_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout112_A hold176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3626_ _3631_/CLK _3626_/D _3117_/Y vssd1 vssd1 vccd1 vccd1 _3626_/Q sky130_fd_sc_hd__dfrtp_4
X_3557_ _3559_/CLK _3557_/D _3051_/Y vssd1 vssd1 vccd1 vccd1 _3557_/Q sky130_fd_sc_hd__dfrtp_1
X_2508_ _2508_/A _2508_/B _2508_/C vssd1 vssd1 vccd1 vccd1 _2568_/D sky130_fd_sc_hd__and3_2
X_3488_ _3488_/CLK _3488_/D _2982_/Y vssd1 vssd1 vccd1 vccd1 _3488_/Q sky130_fd_sc_hd__dfrtp_1
X_2439_ _2439_/A _2584_/C vssd1 vssd1 vccd1 vccd1 _2508_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_66_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2799__A1 _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1810_ _1810_/A vssd1 vssd1 vccd1 vccd1 _1810_/Y sky130_fd_sc_hd__inv_2
X_2790_ _2810_/A1 hold337/X _2793_/S vssd1 vssd1 vccd1 vccd1 _2790_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1741_ _1741_/A _1741_/B _1741_/C _1741_/D vssd1 vssd1 vccd1 vccd1 _1741_/Y sky130_fd_sc_hd__nor4_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold307 _3251_/Q vssd1 vssd1 vccd1 vccd1 hold307/X sky130_fd_sc_hd__dlygate4sd3_1
X_1672_ _2397_/A _3610_/Q _1675_/S vssd1 vssd1 vccd1 vccd1 _1672_/X sky130_fd_sc_hd__mux2_1
Xhold329 _3292_/Q vssd1 vssd1 vccd1 vccd1 hold329/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 _2781_/X vssd1 vssd1 vccd1 vccd1 _3302_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3411_ _3582_/CLK _3411_/D vssd1 vssd1 vccd1 vccd1 _3411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3342_ _3609_/CLK _3342_/D _2917_/Y vssd1 vssd1 vccd1 vccd1 _3342_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1614__A _2287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _3325_/CLK _3273_/D vssd1 vssd1 vccd1 vccd1 _3273_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1029 _2276_/Y vssd1 vssd1 vccd1 vccd1 _3465_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1007 _1794_/X vssd1 vssd1 vccd1 vccd1 _3439_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 _3438_/Q vssd1 vssd1 vccd1 vccd1 _1808_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ _3491_/Q _2224_/B vssd1 vssd1 vccd1 vccd1 _2243_/C sky130_fd_sc_hd__or2_1
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2155_ _2129_/A _3496_/Q _2152_/Y _2130_/B vssd1 vssd1 vccd1 vccd1 _2155_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_88_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2086_ _2121_/A _3544_/Q _2056_/A _2084_/Y vssd1 vssd1 vccd1 vccd1 _2086_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_48_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2650__A0 _2339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2988_ _3105_/A vssd1 vssd1 vccd1 vccd1 _2988_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_56_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1939_ _1926_/Y _1933_/Y _1938_/X _1933_/B _2350_/B vssd1 vssd1 vccd1 vccd1 _1939_/X
+ sky130_fd_sc_hd__a32o_1
X_3609_ _3609_/CLK _3609_/D _3100_/Y vssd1 vssd1 vccd1 vccd1 _3609_/Q sky130_fd_sc_hd__dfrtp_1
Xhold830 _3550_/Q vssd1 vssd1 vccd1 vccd1 hold830/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 _2237_/Y vssd1 vssd1 vccd1 vccd1 _2238_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold852 _1700_/Y vssd1 vssd1 vccd1 vccd1 _3466_/D sky130_fd_sc_hd__clkbuf_2
Xhold863 _3441_/Q vssd1 vssd1 vccd1 vccd1 _1808_/A sky130_fd_sc_hd__buf_1
Xhold896 _2284_/X vssd1 vssd1 vccd1 vccd1 _3461_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 _3466_/Q vssd1 vssd1 vccd1 vccd1 _2258_/S sky130_fd_sc_hd__buf_1
Xhold874 _3549_/Q vssd1 vssd1 vccd1 vccd1 hold874/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2339__B _2339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2880__A0 _2111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1683__A1 hold44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2632__A0 _2342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2911_ _2079_/A hold598/X _2914_/S vssd1 vssd1 vccd1 vccd1 _2911_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2842_ _2338_/B hold746/X _2843_/S vssd1 vssd1 vccd1 vccd1 _2842_/X sky130_fd_sc_hd__mux2_1
X_2773_ _2813_/A1 hold461/X _2773_/S vssd1 vssd1 vccd1 vccd1 _2773_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1724_ _1847_/A _3453_/Q _1722_/X _1723_/X vssd1 vssd1 vccd1 vccd1 _1743_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_13_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1609__A _1609_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold104 _1632_/X vssd1 vssd1 vccd1 vccd1 _3636_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 input29/X vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold115 _1658_/B vssd1 vssd1 vccd1 vccd1 _1669_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 _3198_/Q vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 _2592_/X vssd1 vssd1 vccd1 vccd1 _3137_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1655_ hold288/X _2395_/A hold60/X vssd1 vssd1 vccd1 vccd1 _3616_/D sky130_fd_sc_hd__mux2_1
Xhold148 _3299_/Q vssd1 vssd1 vccd1 vccd1 hold148/X sky130_fd_sc_hd__dlygate4sd3_1
X_1586_ _1838_/B vssd1 vssd1 vccd1 vccd1 _1881_/A sky130_fd_sc_hd__inv_2
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2699__A0 _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ _3325_/CLK _3325_/D vssd1 vssd1 vccd1 vccd1 _3325_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _3331_/CLK _3256_/D vssd1 vssd1 vccd1 vccd1 _3256_/Q sky130_fd_sc_hd__dfxtp_1
X_2207_ _2207_/A _2207_/B vssd1 vssd1 vccd1 vccd1 _2216_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3187_ _3436_/CLK _3187_/D vssd1 vssd1 vccd1 vccd1 _3187_/Q sky130_fd_sc_hd__dfxtp_1
X_2138_ _2134_/B _2134_/C _2136_/C _2134_/A vssd1 vssd1 vccd1 vccd1 _2139_/B sky130_fd_sc_hd__a31o_1
X_2069_ _2121_/A _2069_/B vssd1 vssd1 vccd1 vccd1 _2069_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2623__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold671 _2886_/X vssd1 vssd1 vccd1 vccd1 _3410_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold660 _3368_/Q vssd1 vssd1 vccd1 vccd1 hold660/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 _2645_/X vssd1 vssd1 vccd1 vccd1 _3182_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 _3163_/Q vssd1 vssd1 vccd1 vccd1 hold682/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2318__B1_N _2039_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2862__A0 _2075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1665__A1 _2396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2614__A0 _2111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3110_ _3114_/A vssd1 vssd1 vccd1 vccd1 _3110_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3041_ _3073_/A vssd1 vssd1 vccd1 vccd1 _3041_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2528__S0 _1911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2853__A0 _2339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1656__A1 _2585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1611__B hold65/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2605__A0 _2079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2825_ hold546/X _2342_/B _2833_/S vssd1 vssd1 vccd1 vccd1 _2825_/X sky130_fd_sc_hd__mux2_1
X_2756_ hold189/X _2806_/A1 _2763_/S vssd1 vssd1 vccd1 vccd1 _2756_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1707_ _1707_/A _1707_/B vssd1 vssd1 vccd1 vccd1 _1707_/Y sky130_fd_sc_hd__nand2_1
X_2687_ _2807_/A1 hold229/X _2693_/S vssd1 vssd1 vccd1 vccd1 _2687_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1638_ hold90/X hold52/X hold8/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__mux2_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1569_ _3620_/Q vssd1 vssd1 vccd1 vccd1 _1569_/Y sky130_fd_sc_hd__inv_2
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3308_ _3318_/CLK _3308_/D vssd1 vssd1 vccd1 vccd1 _3308_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2519__S0 _2554_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ _3513_/CLK _3239_/D vssd1 vssd1 vccd1 vccd1 _3239_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout98 _2224_/B vssd1 vssd1 vccd1 vccd1 _1590_/A sky130_fd_sc_hd__buf_8
XFILLER_0_64_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout87 _1911_/C vssd1 vssd1 vccd1 vccd1 _1943_/B sky130_fd_sc_hd__buf_8
Xfanout76 _1745_/Y vssd1 vssd1 vccd1 vccd1 _2383_/C sky130_fd_sc_hd__buf_4
XFILLER_0_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold490 _1939_/X vssd1 vssd1 vccd1 vccd1 _3516_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2835__A0 _2342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1638__A1 hold52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3590_ _3633_/CLK hold53/X _3081_/Y vssd1 vssd1 vccd1 vccd1 _3590_/Q sky130_fd_sc_hd__dfrtp_1
X_2610_ _2342_/B hold676/X _2618_/S vssd1 vssd1 vccd1 vccd1 _2610_/X sky130_fd_sc_hd__mux2_1
X_2541_ _3408_/Q _3399_/Q _3390_/Q _3435_/Q _1943_/B _2550_/S1 vssd1 vssd1 vccd1 vccd1
+ _2541_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2689__S _2693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2472_ _2471_/X _2468_/X _3522_/Q vssd1 vssd1 vccd1 vccd1 _2472_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1972__S1 _2193_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3024_ _3036_/A vssd1 vssd1 vccd1 vccd1 _3024_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_13_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3316_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_18_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2808_ hold140/X _2808_/A1 _2813_/S vssd1 vssd1 vccd1 vccd1 _2808_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_41_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2739_ _2809_/A1 hold422/X _2743_/S vssd1 vssd1 vccd1 vccd1 _2739_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2348__A2 _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1972_ _3249_/Q _3321_/Q _3312_/Q _3303_/Q _1590_/A _2193_/A1 vssd1 vssd1 vccd1 vccd1
+ _1972_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_28_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3642_ _3642_/CLK hold97/X _3133_/Y vssd1 vssd1 vccd1 vccd1 _3642_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_70_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3573_ _3576_/CLK _3573_/D _3067_/Y vssd1 vssd1 vccd1 vccd1 _3573_/Q sky130_fd_sc_hd__dfrtp_1
X_2524_ hold78/A _2568_/B _2417_/B _3378_/Q _2523_/X vssd1 vssd1 vccd1 vccd1 _2524_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2455_ _2506_/S _2454_/X _2447_/X vssd1 vssd1 vccd1 vccd1 _2455_/X sky130_fd_sc_hd__a21o_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_2386_ hold74/A _3380_/Q _3377_/Q hold79/A vssd1 vssd1 vccd1 vccd1 _2386_/X sky130_fd_sc_hd__a22o_1
X_3007_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3007_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_2_1__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2792__S _2793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ _2367_/B _1889_/Y _2231_/A vssd1 vssd1 vccd1 vccd1 _2241_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__3652__A _3659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2171_ _2794_/A _2175_/A vssd1 vssd1 vccd1 vccd1 _2228_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__3099__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1955_ _3346_/Q _2379_/S vssd1 vssd1 vccd1 vccd1 _1955_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1886_ _1602_/Y _1603_/Y _1813_/A _1745_/B vssd1 vssd1 vccd1 vccd1 _2915_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_43_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3625_ _3629_/CLK _3625_/D _3116_/Y vssd1 vssd1 vccd1 vccd1 _3625_/Q sky130_fd_sc_hd__dfrtp_4
X_3556_ _3559_/CLK _3556_/D _3050_/Y vssd1 vssd1 vccd1 vccd1 _3556_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout105_A hold86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2507_ hold59/A _2507_/B _2507_/C vssd1 vssd1 vccd1 vccd1 _2508_/C sky130_fd_sc_hd__and3_1
X_3487_ _3488_/CLK _3487_/D _2981_/Y vssd1 vssd1 vccd1 vccd1 _3487_/Q sky130_fd_sc_hd__dfrtp_1
X_2438_ _3612_/Q _2439_/A _2406_/X vssd1 vssd1 vccd1 vccd1 _2438_/X sky130_fd_sc_hd__a21o_1
X_2369_ hold70/X hold90/X hold80/X vssd1 vssd1 vccd1 vccd1 _2370_/A sky130_fd_sc_hd__or3_2
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2787__S _2793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1740_ _1853_/A _2580_/A _1715_/X _1716_/X _1717_/X vssd1 vssd1 vccd1 vccd1 _1740_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_25_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold308 _2725_/X vssd1 vssd1 vccd1 vccd1 _3251_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1671_ _2585_/B _1671_/B vssd1 vssd1 vccd1 vccd1 _1671_/Y sky130_fd_sc_hd__nand2_1
Xhold319 _3301_/Q vssd1 vssd1 vccd1 vccd1 hold319/X sky130_fd_sc_hd__dlygate4sd3_1
X_3410_ _3423_/CLK _3410_/D vssd1 vssd1 vccd1 vccd1 _3410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3341_ _3580_/CLK _3341_/D _1606_/Y vssd1 vssd1 vccd1 vccd1 _3341_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _3318_/CLK _3272_/D vssd1 vssd1 vccd1 vccd1 _3272_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1008 _3463_/Q vssd1 vssd1 vccd1 vccd1 _2273_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1019 _2374_/X vssd1 vssd1 vccd1 vccd1 _3438_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2022__S0 _2044_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ _3491_/Q _2224_/B vssd1 vssd1 vccd1 vccd1 _2243_/B sky130_fd_sc_hd__nand2_1
X_2154_ _2130_/A _3347_/Q _2156_/A _2152_/Y hold989/X vssd1 vssd1 vccd1 vccd1 _2154_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_23_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2085_ _3544_/Q _2089_/B vssd1 vssd1 vccd1 vccd1 _2085_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2987_ _3105_/A vssd1 vssd1 vccd1 vccd1 _2987_/Y sky130_fd_sc_hd__inv_2
X_1938_ _3515_/Q _1938_/B vssd1 vssd1 vccd1 vccd1 _1938_/X sky130_fd_sc_hd__or2_1
X_1869_ _3534_/Q _3533_/Q _1843_/B _1845_/A vssd1 vssd1 vccd1 vccd1 _1869_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3608_ _3609_/CLK _3608_/D _3099_/Y vssd1 vssd1 vccd1 vccd1 _3608_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold820 _3506_/Q vssd1 vssd1 vccd1 vccd1 hold820/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 _3469_/Q vssd1 vssd1 vccd1 vccd1 hold853/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold831 _1827_/X vssd1 vssd1 vccd1 vccd1 _3549_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 _2384_/X vssd1 vssd1 vccd1 vccd1 _3441_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 _2238_/Y vssd1 vssd1 vccd1 vccd1 _3479_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3539_ _3539_/CLK _3539_/D _3033_/Y vssd1 vssd1 vccd1 vccd1 _3539_/Q sky130_fd_sc_hd__dfrtp_1
Xhold897 _3577_/Q vssd1 vssd1 vccd1 vccd1 _1701_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 _3503_/Q vssd1 vssd1 vccd1 vccd1 _2125_/A sky130_fd_sc_hd__buf_1
Xhold886 _3580_/Q vssd1 vssd1 vccd1 vccd1 hold886/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2013__S0 _1590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2910_ _2111_/B hold776/X _2914_/S vssd1 vssd1 vccd1 vccd1 _2910_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2841_ _2075_/B hold684/X _2843_/S vssd1 vssd1 vccd1 vccd1 _2841_/X sky130_fd_sc_hd__mux2_1
X_2772_ _2812_/A1 hold292/X _2773_/S vssd1 vssd1 vccd1 vccd1 _2772_/X sky130_fd_sc_hd__mux2_1
X_1723_ _3457_/Q _1859_/A vssd1 vssd1 vccd1 vccd1 _1723_/X sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_38_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3582_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1609__B _1609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold105 _3619_/Q vssd1 vssd1 vccd1 vccd1 hold105/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold116 _2441_/A vssd1 vssd1 vccd1 vccd1 _1671_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 _1672_/X vssd1 vssd1 vccd1 vccd1 _3610_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _2778_/X vssd1 vssd1 vccd1 vccd1 _3299_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _3227_/Q vssd1 vssd1 vccd1 vccd1 hold138/X sky130_fd_sc_hd__dlygate4sd3_1
X_1654_ _1571_/A _2396_/A hold60/X vssd1 vssd1 vccd1 vccd1 _3617_/D sky130_fd_sc_hd__mux2_1
X_1585_ _1838_/A vssd1 vssd1 vccd1 vccd1 _1879_/A sky130_fd_sc_hd__inv_2
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3324_ _3328_/CLK _3324_/D vssd1 vssd1 vccd1 vccd1 _3324_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3330_/CLK _3255_/D vssd1 vssd1 vccd1 vccd1 _3255_/Q sky130_fd_sc_hd__dfxtp_1
X_2206_ _3483_/Q _2218_/B vssd1 vssd1 vccd1 vccd1 _2207_/B sky130_fd_sc_hd__nand2_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _3435_/CLK _3186_/D vssd1 vssd1 vccd1 vccd1 _3186_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2871__A1 _2079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2137_ _2125_/A _2139_/A _2136_/X vssd1 vssd1 vccd1 vccd1 _2137_/X sky130_fd_sc_hd__a21o_1
X_2068_ _2080_/A _2068_/B vssd1 vssd1 vccd1 vccd1 _2076_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_88_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2890__S _2894_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold650 _3171_/Q vssd1 vssd1 vccd1 vccd1 hold650/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 _2845_/X vssd1 vssd1 vccd1 vccd1 _3368_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 _3409_/Q vssd1 vssd1 vccd1 vccd1 hold672/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 _3174_/Q vssd1 vssd1 vccd1 vccd1 hold694/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 _2623_/X vssd1 vssd1 vccd1 vccd1 _3163_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout85_A _1942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output66_A _2562_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3040_ _3073_/A vssd1 vssd1 vccd1 vccd1 _3040_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2528__S1 _2550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1611__C input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2824_ _2895_/C _2824_/B _2905_/B vssd1 vssd1 vccd1 vccd1 _2833_/S sky130_fd_sc_hd__and3b_4
XFILLER_0_14_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2755_ hold309/X _2805_/A1 _2763_/S vssd1 vssd1 vccd1 vccd1 _2755_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1706_ _1703_/B hold903/X _3466_/D vssd1 vssd1 vccd1 vccd1 _1706_/Y sky130_fd_sc_hd__a21oi_1
X_2686_ _2806_/A1 hold181/X _2693_/S vssd1 vssd1 vccd1 vccd1 _2686_/X sky130_fd_sc_hd__mux2_1
X_1637_ hold70/X hold44/X hold8/X vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3307_ _3316_/CLK _3307_/D vssd1 vssd1 vccd1 vccd1 _3307_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1568_ hold87/X vssd1 vssd1 vccd1 vccd1 _1568_/Y sky130_fd_sc_hd__inv_2
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2519__S1 _1911_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3238_ _3328_/CLK _3238_/D vssd1 vssd1 vccd1 vccd1 _3238_/Q sky130_fd_sc_hd__dfxtp_1
X_3169_ _3433_/CLK _3169_/D vssd1 vssd1 vccd1 vccd1 _3169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout99 hold501/X vssd1 vssd1 vccd1 vccd1 _2224_/B sky130_fd_sc_hd__buf_4
XFILLER_0_64_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout88 _1911_/C vssd1 vssd1 vccd1 vccd1 _2554_/S0 sky130_fd_sc_hd__buf_6
XFILLER_0_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2780__A0 _2810_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold480 _1949_/X vssd1 vssd1 vccd1 vccd1 _3514_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 _3521_/Q vssd1 vssd1 vccd1 vccd1 _1911_/A sky130_fd_sc_hd__buf_1
XFILLER_0_87_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3655__A _3659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2540_ _2511_/Y _2538_/X _2539_/X _2511_/B hold62/A vssd1 vssd1 vccd1 vccd1 _2540_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__2771__A0 _2811_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2471_ _2470_/X _2469_/X _3521_/Q vssd1 vssd1 vccd1 vccd1 _2471_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3023_ _3036_/A vssd1 vssd1 vccd1 vccd1 _3023_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2826__A1 _2097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2807_ hold248/X _2807_/A1 _2813_/S vssd1 vssd1 vccd1 vccd1 _2807_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2738_ _2808_/A1 hold150/X _2743_/S vssd1 vssd1 vccd1 vccd1 _2738_/X sky130_fd_sc_hd__mux2_1
X_2669_ _2810_/A1 hold323/X _2672_/S vssd1 vssd1 vccd1 vccd1 _2669_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2817__A1 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2428__S0 _1943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2753__A0 _2813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2808__A1 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1971_ _3294_/Q _3285_/Q _3276_/Q _3267_/Q _1590_/A _2193_/A1 vssd1 vssd1 vccd1 vccd1
+ _1971_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_55_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3641_ _3642_/CLK _3641_/D _3132_/Y vssd1 vssd1 vccd1 vccd1 _3641_/Q sky130_fd_sc_hd__dfrtp_1
X_3572_ _3576_/CLK _3572_/D _3066_/Y vssd1 vssd1 vccd1 vccd1 _3572_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2523_ _3590_/Q hold67/A vssd1 vssd1 vccd1 vccd1 _2523_/X sky130_fd_sc_hd__or2_1
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2454_ _2453_/X _2450_/X _3522_/Q vssd1 vssd1 vccd1 vccd1 _2454_/X sky130_fd_sc_hd__mux2_1
X_2385_ _1811_/A _1795_/B _2381_/B _1775_/Y _1815_/B vssd1 vssd1 vccd1 vccd1 _2385_/X
+ sky130_fd_sc_hd__a32o_1
Xinput1 uart_rx vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3006_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3006_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2735__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2726__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2170_ _2794_/B _2179_/A _3491_/Q vssd1 vssd1 vccd1 vccd1 _2175_/A sky130_fd_sc_hd__and3_1
XFILLER_0_73_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1954_ _2366_/A _2366_/B vssd1 vssd1 vccd1 vccd1 _2379_/S sky130_fd_sc_hd__nand2_1
XFILLER_0_83_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1885_ _1835_/A _1560_/Y _1885_/S vssd1 vssd1 vccd1 vccd1 _3527_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_3_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3624_ _3629_/CLK _3624_/D _3115_/Y vssd1 vssd1 vccd1 vccd1 _3624_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__2717__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3555_ _3563_/CLK _3555_/D _3049_/Y vssd1 vssd1 vccd1 vccd1 _3555_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2193__A1 _2193_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3486_ _3610_/CLK _3486_/D _2980_/Y vssd1 vssd1 vccd1 vccd1 _3486_/Q sky130_fd_sc_hd__dfrtp_1
X_2506_ _2498_/X _2505_/X _2506_/S vssd1 vssd1 vccd1 vccd1 _2506_/X sky130_fd_sc_hd__mux2_1
X_2437_ _3616_/Q _1645_/Y _2571_/B vssd1 vssd1 vccd1 vccd1 _2437_/X sky130_fd_sc_hd__a21o_1
X_2368_ _2052_/S _2366_/X _2367_/X _1600_/Y vssd1 vssd1 vccd1 vccd1 _2368_/Y sky130_fd_sc_hd__o22ai_1
X_2299_ hold98/X hold49/X hold30/X vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__mux2_1
XANTENNA__2893__S _2894_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2708__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1670_ _2441_/A vssd1 vssd1 vccd1 vccd1 _2476_/B sky130_fd_sc_hd__inv_2
XFILLER_0_13_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold309 _3278_/Q vssd1 vssd1 vccd1 vccd1 hold309/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3340_ _3433_/CLK _3340_/D vssd1 vssd1 vccd1 vccd1 _3340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3305_/CLK _3271_/D vssd1 vssd1 vccd1 vccd1 _3271_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1009 _2279_/Y vssd1 vssd1 vccd1 vccd1 _2280_/C sky130_fd_sc_hd__dlygate4sd3_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2022__S1 _2044_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2222_ _2222_/A _2222_/B vssd1 vssd1 vccd1 vccd1 _2226_/A sky130_fd_sc_hd__xnor2_1
X_2153_ _2147_/Y _2161_/S _1589_/A vssd1 vssd1 vccd1 vccd1 _2153_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2084_ _2121_/A _2084_/B vssd1 vssd1 vccd1 vccd1 _2084_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_75_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2986_ _3105_/A vssd1 vssd1 vccd1 vccd1 _2986_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_56_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1937_ _1930_/X _1936_/Y _1928_/A _1933_/B vssd1 vssd1 vccd1 vccd1 _3517_/D sky130_fd_sc_hd__a2bb2o_1
X_1868_ _1867_/Y _1865_/B _1584_/A _1560_/Y vssd1 vssd1 vccd1 vccd1 _3536_/D sky130_fd_sc_hd__a2bb2o_1
X_3607_ _3609_/CLK _3607_/D _3098_/Y vssd1 vssd1 vccd1 vccd1 _3607_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2888__S _2894_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold821 _2042_/X vssd1 vssd1 vccd1 vccd1 _3506_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold810 _3512_/Q vssd1 vssd1 vccd1 vccd1 hold810/X sky130_fd_sc_hd__dlygate4sd3_1
X_3538_ _3540_/CLK _3538_/D _3032_/Y vssd1 vssd1 vccd1 vccd1 _3538_/Q sky130_fd_sc_hd__dfrtp_1
Xhold843 _3472_/Q vssd1 vssd1 vccd1 vccd1 hold843/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold854 _2256_/X vssd1 vssd1 vccd1 vccd1 _3470_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1799_ _1778_/A _1824_/A _1803_/B _1799_/D vssd1 vssd1 vccd1 vccd1 _1799_/X sky130_fd_sc_hd__and4b_1
Xhold832 _3507_/Q vssd1 vssd1 vccd1 vccd1 hold832/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 _3471_/Q vssd1 vssd1 vccd1 vccd1 hold865/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 _1701_/Y vssd1 vssd1 vccd1 vccd1 hold898/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 _2137_/X vssd1 vssd1 vccd1 vccd1 _3503_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 _2916_/X vssd1 vssd1 vccd1 vccd1 _3580_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3469_ _3583_/CLK _3469_/D _2963_/Y vssd1 vssd1 vccd1 vccd1 _3469_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2013__S1 _2222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_8_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3330_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1967__S _2053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2840_ _2079_/A hold638/X _2843_/S vssd1 vssd1 vccd1 vccd1 _2840_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3658__A _3659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2771_ _2811_/A1 hold434/X _2773_/S vssd1 vssd1 vccd1 vccd1 _2771_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1722_ _1582_/Y _3459_/Q hold204/X _1879_/A vssd1 vssd1 vccd1 vccd1 _1722_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_5_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1609__C _1907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold117 _1671_/Y vssd1 vssd1 vccd1 vccd1 _1675_/S sky130_fd_sc_hd__clkbuf_2
X_1653_ _1570_/A _2397_/A hold60/X vssd1 vssd1 vccd1 vccd1 _3618_/D sky130_fd_sc_hd__mux2_1
Xhold106 _3628_/Q vssd1 vssd1 vccd1 vccd1 _2383_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold139 _2698_/X vssd1 vssd1 vccd1 vccd1 _3227_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 _3254_/Q vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
X_1584_ _1584_/A vssd1 vssd1 vccd1 vccd1 _1847_/A sky130_fd_sc_hd__inv_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1625__B _1625_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3323_ _3325_/CLK _3323_/D vssd1 vssd1 vccd1 vccd1 _3323_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ _3328_/CLK _3254_/D vssd1 vssd1 vccd1 vccd1 _3254_/Q sky130_fd_sc_hd__dfxtp_1
X_2205_ _2205_/A _2211_/B vssd1 vssd1 vccd1 vccd1 _2218_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_28_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ _3435_/CLK _3185_/D vssd1 vssd1 vccd1 vccd1 _3185_/Q sky130_fd_sc_hd__dfxtp_1
X_2136_ _2125_/A _3346_/Q _2136_/C _2136_/D vssd1 vssd1 vccd1 vccd1 _2136_/X sky130_fd_sc_hd__and4b_1
X_2067_ _2082_/A _2067_/B _2082_/B vssd1 vssd1 vccd1 vccd1 _2067_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_88_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2969_ _3073_/A vssd1 vssd1 vccd1 vccd1 _2969_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold640 _3183_/Q vssd1 vssd1 vccd1 vccd1 hold640/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 _2633_/X vssd1 vssd1 vccd1 vccd1 _3171_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 _3192_/Q vssd1 vssd1 vccd1 vccd1 hold662/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 _2636_/X vssd1 vssd1 vccd1 vccd1 _3174_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 _3365_/Q vssd1 vssd1 vccd1 vccd1 hold684/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 _2884_/X vssd1 vssd1 vccd1 vccd1 _3409_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2302__A1 hold33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1611__D input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2823_ hold522/X _2339_/B _2823_/S vssd1 vssd1 vccd1 vccd1 _2823_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2754_ _2794_/C _2794_/A _2794_/B vssd1 vssd1 vccd1 vccd1 _2763_/S sky130_fd_sc_hd__nor3b_4
XFILLER_0_60_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1705_ _1705_/A _1705_/B vssd1 vssd1 vccd1 vccd1 _1705_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2685_ _2805_/A1 hold242/X _2693_/S vssd1 vssd1 vccd1 vccd1 _2685_/X sky130_fd_sc_hd__mux2_1
X_1636_ hold54/X hold49/X hold8/X vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1567_ _2121_/A vssd1 vssd1 vccd1 vccd1 _2071_/A sky130_fd_sc_hd__inv_2
X_3306_ _3319_/CLK _3306_/D vssd1 vssd1 vccd1 vccd1 _3306_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _3331_/CLK _3237_/D vssd1 vssd1 vccd1 vccd1 _3237_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3168_ _3435_/CLK _3168_/D vssd1 vssd1 vccd1 vccd1 _3168_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2186__B _2200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2119_ _2114_/Y _2116_/X _2118_/X _1772_/B _1605_/Y vssd1 vssd1 vccd1 vccd1 _2119_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3099_ _3126_/A vssd1 vssd1 vccd1 vccd1 _3099_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_76_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout89 hold483/X vssd1 vssd1 vccd1 vccd1 _1911_/C sky130_fd_sc_hd__clkbuf_8
Xfanout78 _2067_/Y vssd1 vssd1 vccd1 vccd1 _2079_/A sky130_fd_sc_hd__buf_4
XFILLER_0_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold470 _3486_/Q vssd1 vssd1 vccd1 vccd1 _2211_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold481 _3581_/Q vssd1 vssd1 vccd1 vccd1 _2586_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 _3522_/Q vssd1 vssd1 vccd1 vccd1 _1912_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2470_ _3172_/Q _3421_/Q _3412_/Q _3154_/Q _2554_/S0 _1911_/B vssd1 vssd1 vccd1 vccd1
+ _2470_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2287__A _2287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3022_ _3036_/A vssd1 vssd1 vccd1 vccd1 _3022_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_58_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout128_A _3131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2806_ hold183/X _2806_/A1 _2813_/S vssd1 vssd1 vccd1 vccd1 _2806_/X sky130_fd_sc_hd__mux2_1
X_2737_ _2807_/A1 hold231/X _2743_/S vssd1 vssd1 vccd1 vccd1 _2737_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_22_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3636_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2762__A1 _2812_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2668_ _2809_/A1 hold358/X _2672_/S vssd1 vssd1 vccd1 vccd1 _2668_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2896__S _2904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1619_ _3642_/Q hold86/X _1623_/S vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__mux2_1
X_2599_ _2824_/B _2905_/B _2905_/C vssd1 vssd1 vccd1 vccd1 _2608_/S sky130_fd_sc_hd__or3b_4
XFILLER_0_69_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2428__S1 _1942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1970_ _1968_/X _1969_/X _2045_/S vssd1 vssd1 vccd1 vccd1 _1970_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2570__A _2583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3640_ _3642_/CLK _3640_/D _3131_/Y vssd1 vssd1 vccd1 vccd1 _3640_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3571_ _3571_/CLK _3571_/D _3065_/Y vssd1 vssd1 vccd1 vccd1 _3571_/Q sky130_fd_sc_hd__dfstp_1
X_2522_ _2583_/B _2514_/X _2521_/X _2506_/S vssd1 vssd1 vccd1 vccd1 _2522_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_87_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2453_ _2452_/X _2451_/X _2551_/S vssd1 vssd1 vccd1 vccd1 _2453_/X sky130_fd_sc_hd__mux2_1
X_2384_ _1808_/A _1772_/B _2383_/X vssd1 vssd1 vccd1 vccd1 _2384_/X sky130_fd_sc_hd__a21o_1
Xinput2 wb_rst_i vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_1
X_3005_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3005_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2671__A0 _2812_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output41_A _2435_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1953_ _2130_/A _2156_/A vssd1 vssd1 vccd1 vccd1 _2366_/B sky130_fd_sc_hd__and2_2
X_1884_ _1835_/A _1881_/B _1883_/X _1883_/A _1560_/Y vssd1 vssd1 vccd1 vccd1 _1884_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__2504__S _2551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3623_ _3623_/CLK hold50/X _3114_/Y vssd1 vssd1 vccd1 vccd1 _3623_/Q sky130_fd_sc_hd__dfrtp_1
X_3554_ _3559_/CLK _3554_/D _3048_/Y vssd1 vssd1 vccd1 vccd1 _3554_/Q sky130_fd_sc_hd__dfrtp_1
X_3485_ _3609_/CLK _3485_/D _2979_/Y vssd1 vssd1 vccd1 vccd1 _3485_/Q sky130_fd_sc_hd__dfrtp_1
X_2505_ _2501_/X _2504_/X _3522_/Q vssd1 vssd1 vccd1 vccd1 _2505_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2193__A2 _2224_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2436_ _3639_/Q _2511_/A _2511_/B vssd1 vssd1 vccd1 vccd1 _2436_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2367_ _2367_/A _2367_/B _2367_/C vssd1 vssd1 vccd1 vccd1 _2367_/X sky130_fd_sc_hd__or3_1
X_2298_ _3453_/Q hold14/X hold30/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__mux2_1
XANTENNA__2653__A0 _2097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2500__S0 _2554_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2644__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3270_ _3319_/CLK _3270_/D vssd1 vssd1 vccd1 vccd1 _3270_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _3492_/Q _3491_/Q vssd1 vssd1 vccd1 vccd1 _2222_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_84_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1686__A1 hold86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2883__A0 _2338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2152_ _2161_/S vssd1 vssd1 vccd1 vccd1 _2152_/Y sky130_fd_sc_hd__inv_2
X_2083_ _3545_/Q _2089_/B vssd1 vssd1 vccd1 vccd1 _2084_/B sky130_fd_sc_hd__nand2_1
XANTENNA__1911__B _1911_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2635__A0 _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2985_ _3105_/A vssd1 vssd1 vccd1 vccd1 _2985_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_71_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1936_ _1930_/A _1930_/B _1933_/Y vssd1 vssd1 vccd1 vccd1 _1936_/Y sky130_fd_sc_hd__o21ai_1
X_1867_ _1584_/A _1846_/A _1835_/A vssd1 vssd1 vccd1 vccd1 _1867_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold800 _3385_/Q vssd1 vssd1 vccd1 vccd1 hold800/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout110_A hold120/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1798_ _1604_/Y _1799_/D _1803_/B vssd1 vssd1 vccd1 vccd1 _1802_/A sky130_fd_sc_hd__o21ai_1
Xhold811 _1978_/X vssd1 vssd1 vccd1 vccd1 _3512_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3606_ _3614_/CLK _3606_/D _3097_/Y vssd1 vssd1 vccd1 vccd1 _3606_/Q sky130_fd_sc_hd__dfrtp_1
X_3537_ _3539_/CLK _3537_/D _3031_/Y vssd1 vssd1 vccd1 vccd1 _3537_/Q sky130_fd_sc_hd__dfrtp_1
Xhold844 _2253_/X vssd1 vssd1 vccd1 vccd1 _3473_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 _3551_/Q vssd1 vssd1 vccd1 vccd1 hold855/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 _2031_/X vssd1 vssd1 vccd1 vccd1 _3507_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold822 _3513_/Q vssd1 vssd1 vccd1 vccd1 hold822/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 _3543_/Q vssd1 vssd1 vccd1 vccd1 hold888/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold866 _2255_/X vssd1 vssd1 vccd1 vccd1 _3471_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold877 _3545_/Q vssd1 vssd1 vccd1 vccd1 hold877/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 _1702_/Y vssd1 vssd1 vccd1 vccd1 _3577_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3468_ _3583_/CLK _3468_/D _2962_/Y vssd1 vssd1 vccd1 vccd1 _3468_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2549__S0 _1911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3399_ _3435_/CLK _3399_/D vssd1 vssd1 vccd1 vccd1 _3399_/Q sky130_fd_sc_hd__dfxtp_1
X_2419_ _2419_/A _2419_/B vssd1 vssd1 vccd1 vccd1 _2584_/C sky130_fd_sc_hd__and2_1
XANTENNA__2626__A0 _2079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2617__A0 _2338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2770_ _2810_/A1 hold329/X _2773_/S vssd1 vssd1 vccd1 vccd1 _2770_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1721_ _1845_/A hold98/X vssd1 vssd1 vccd1 vccd1 _1721_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_80_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold107 _1640_/X vssd1 vssd1 vccd1 vccd1 _3628_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1652_ hold105/X hold86/X hold60/X vssd1 vssd1 vccd1 vccd1 _3619_/D sky130_fd_sc_hd__mux2_1
Xhold118 _1675_/X vssd1 vssd1 vccd1 vccd1 _3607_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 _2728_/X vssd1 vssd1 vccd1 vccd1 _3254_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1583_ _1583_/A vssd1 vssd1 vccd1 vccd1 _1851_/A sky130_fd_sc_hd__inv_2
X_3322_ _3483_/CLK _3322_/D vssd1 vssd1 vccd1 vccd1 _3322_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _3330_/CLK _3253_/D vssd1 vssd1 vccd1 vccd1 _3253_/Q sky130_fd_sc_hd__dfxtp_1
X_2204_ _2205_/A _2211_/B vssd1 vssd1 vccd1 vccd1 _2207_/A sky130_fd_sc_hd__nand2_1
X_3184_ _3435_/CLK _3184_/D vssd1 vssd1 vccd1 vccd1 _3184_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_47_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3435_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2856__A0 _2342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2135_ _2052_/S _2136_/D _2136_/C vssd1 vssd1 vccd1 vccd1 _2139_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2608__A0 _2339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2066_ _2060_/Y _2062_/B _2071_/B _2069_/B _2121_/A _2080_/A vssd1 vssd1 vccd1 vccd1
+ _2082_/B sky130_fd_sc_hd__mux4_2
XFILLER_0_88_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2968_ _3073_/A vssd1 vssd1 vccd1 vccd1 _2968_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2899__S _2904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1919_ _1911_/B _1917_/X _1918_/Y _1910_/B vssd1 vssd1 vccd1 vccd1 _1919_/X sky130_fd_sc_hd__o22a_1
X_2899_ hold544/X _2104_/X _2904_/S vssd1 vssd1 vccd1 vccd1 _2899_/X sky130_fd_sc_hd__mux2_1
Xhold630 _3403_/Q vssd1 vssd1 vccd1 vccd1 hold630/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold663 _2656_/X vssd1 vssd1 vccd1 vccd1 _3192_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold641 _2646_/X vssd1 vssd1 vccd1 vccd1 _3183_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 _3411_/Q vssd1 vssd1 vccd1 vccd1 hold652/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 _3156_/Q vssd1 vssd1 vccd1 vccd1 hold696/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 _3372_/Q vssd1 vssd1 vccd1 vccd1 hold674/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 _2841_/X vssd1 vssd1 vccd1 vccd1 _3365_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1978__S _2053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2838__A0 _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2573__A _2583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2822_ hold624/X _2338_/B _2823_/S vssd1 vssd1 vccd1 vccd1 _2822_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2753_ _2813_/A1 hold380/X _2753_/S vssd1 vssd1 vccd1 vccd1 _2753_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1704_ hold908/X _1703_/Y _3466_/D vssd1 vssd1 vccd1 vccd1 _3576_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2684_ _2804_/B _2764_/A vssd1 vssd1 vccd1 vccd1 _2693_/S sky130_fd_sc_hd__or2_4
X_1635_ hold23/X hold14/X hold8/X vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1566_ _3625_/Q vssd1 vssd1 vccd1 vccd1 _1783_/A sky130_fd_sc_hd__inv_2
X_3305_ _3305_/CLK _3305_/D vssd1 vssd1 vccd1 vccd1 _3305_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _3328_/CLK _3236_/D vssd1 vssd1 vccd1 vccd1 _3236_/Q sky130_fd_sc_hd__dfxtp_1
X_3167_ _3436_/CLK _3167_/D vssd1 vssd1 vccd1 vccd1 _3167_/Q sky130_fd_sc_hd__dfxtp_1
X_3098_ _3126_/A vssd1 vssd1 vccd1 vccd1 _3098_/Y sky130_fd_sc_hd__inv_2
X_2118_ hold80/X _2111_/A _2117_/X vssd1 vssd1 vccd1 vccd1 _2118_/X sky130_fd_sc_hd__a21bo_1
X_2049_ _1985_/S _2049_/B vssd1 vssd1 vccd1 vccd1 _2049_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_76_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout68 _2104_/X vssd1 vssd1 vccd1 vccd1 _2105_/B sky130_fd_sc_hd__buf_4
XFILLER_0_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold460 _2723_/X vssd1 vssd1 vccd1 vccd1 _3250_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 _2215_/X vssd1 vssd1 vccd1 vccd1 _3486_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 _3518_/Q vssd1 vssd1 vccd1 vccd1 _1931_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold482 _2586_/Y vssd1 vssd1 vccd1 vccd1 _3581_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2296__A1 hold41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3021_ _3036_/A vssd1 vssd1 vccd1 vccd1 _3021_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2039__A1 _1985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2805_ hold286/X _2805_/A1 _2813_/S vssd1 vssd1 vccd1 vccd1 _2805_/X sky130_fd_sc_hd__mux2_1
X_2736_ _2806_/A1 hold178/X _2743_/S vssd1 vssd1 vccd1 vccd1 _2736_/X sky130_fd_sc_hd__mux2_1
X_2667_ _2808_/A1 hold146/X _2672_/S vssd1 vssd1 vccd1 vccd1 _2667_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1618_ _2393_/A hold96/X vssd1 vssd1 vccd1 vccd1 _1623_/S sky130_fd_sc_hd__nor2_2
XFILLER_0_1_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2598_ _3524_/Q _3523_/Q _2598_/C vssd1 vssd1 vccd1 vccd1 _2905_/C sky130_fd_sc_hd__and3_2
XANTENNA_hold1040_A _3642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3219_ _3331_/CLK _3219_/D vssd1 vssd1 vccd1 vccd1 _3219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold290 _3625_/Q vssd1 vssd1 vccd1 vccd1 _2080_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3570_ _3571_/CLK _3570_/D _3064_/Y vssd1 vssd1 vccd1 vccd1 _3570_/Q sky130_fd_sc_hd__dfstp_1
X_2521_ _2520_/X _2517_/X _3522_/Q vssd1 vssd1 vccd1 vccd1 _2521_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2452_ _3171_/Q _3420_/Q _3411_/Q _3153_/Q _2554_/S0 _1911_/B vssd1 vssd1 vccd1 vccd1
+ _2452_/X sky130_fd_sc_hd__mux4_1
X_2383_ _2383_/A _3438_/Q _2383_/C vssd1 vssd1 vccd1 vccd1 _2383_/X sky130_fd_sc_hd__and3_1
Xinput3 input3/A vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_2
X_3004_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3004_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2680__A1 _2811_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2719_ _2809_/A1 hold420/X _2723_/S vssd1 vssd1 vccd1 vccd1 _2719_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2043__S0 _2044_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1986__S _2052_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2610__S _2618_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1952_ _2130_/B _2129_/A _3496_/Q vssd1 vssd1 vccd1 vccd1 _2156_/A sky130_fd_sc_hd__and3_1
X_1883_ _1883_/A _3527_/Q vssd1 vssd1 vccd1 vccd1 _1883_/X sky130_fd_sc_hd__or2_1
X_3622_ _3631_/CLK _3622_/D _3113_/Y vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3553_ _3559_/CLK _3553_/D _3047_/Y vssd1 vssd1 vccd1 vccd1 _3553_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3484_ _3609_/CLK _3484_/D _2978_/Y vssd1 vssd1 vccd1 vccd1 _3484_/Q sky130_fd_sc_hd__dfrtp_1
X_2504_ _2503_/X _2502_/X _2551_/S vssd1 vssd1 vccd1 vccd1 _2504_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2025__S0 _1590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2435_ _2506_/S _2434_/X _2427_/X vssd1 vssd1 vccd1 vccd1 _2435_/X sky130_fd_sc_hd__a21o_2
X_2366_ _2366_/A _2366_/B _2366_/C vssd1 vssd1 vccd1 vccd1 _2366_/X sky130_fd_sc_hd__and3_1
X_2297_ _3454_/Q hold2/X hold30/A vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__mux2_1
XANTENNA__1660__A _1660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2500__S1 _1911_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2430__S _2551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2341__B1 _2075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1614__C_N _1624_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _2214_/Y _2214_/B _2220_/S vssd1 vssd1 vccd1 vccd1 _2220_/X sky130_fd_sc_hd__mux2_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2576__A _2583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2151_ _2366_/A _2156_/B _2150_/X vssd1 vssd1 vccd1 vccd1 _2161_/S sky130_fd_sc_hd__o21ai_4
X_2082_ _2082_/A _2082_/B vssd1 vssd1 vccd1 vccd1 _2082_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__1911__C _1911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2984_ _3105_/A vssd1 vssd1 vccd1 vccd1 _2984_/Y sky130_fd_sc_hd__inv_2
X_1935_ _1931_/A _1933_/B _1932_/Y _1934_/X vssd1 vssd1 vccd1 vccd1 _1935_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1866_ _1835_/A _1848_/Y _1865_/X _1865_/A _1560_/Y vssd1 vssd1 vccd1 vccd1 _1866_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_31_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3605_ _3633_/CLK hold22/X _3096_/Y vssd1 vssd1 vccd1 vccd1 _3605_/Q sky130_fd_sc_hd__dfrtp_1
Xhold812 _3473_/Q vssd1 vssd1 vccd1 vccd1 hold812/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold801 _2858_/X vssd1 vssd1 vccd1 vccd1 _3385_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1797_ _1797_/A _1797_/B _1803_/A vssd1 vssd1 vccd1 vccd1 _1799_/D sky130_fd_sc_hd__and3_1
X_3536_ _3539_/CLK _3536_/D _3030_/Y vssd1 vssd1 vccd1 vccd1 _3536_/Q sky130_fd_sc_hd__dfrtp_1
Xhold845 _3529_/Q vssd1 vssd1 vccd1 vccd1 _1838_/B sky130_fd_sc_hd__buf_1
Xhold834 _3481_/Q vssd1 vssd1 vccd1 vccd1 _2261_/A sky130_fd_sc_hd__buf_1
XFILLER_0_24_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout103_A hold52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold823 _1967_/X vssd1 vssd1 vccd1 vccd1 _3513_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 _3530_/Q vssd1 vssd1 vccd1 vccd1 _1838_/A sky130_fd_sc_hd__buf_1
Xhold889 _1833_/X vssd1 vssd1 vccd1 vccd1 _3543_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 _1832_/X vssd1 vssd1 vccd1 vccd1 _3544_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 _1826_/X vssd1 vssd1 vccd1 vccd1 _3550_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3467_ _3583_/CLK _3467_/D _2961_/Y vssd1 vssd1 vccd1 vccd1 _3467_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2549__S1 _2550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3398_ _3523_/CLK _3398_/D vssd1 vssd1 vccd1 vccd1 _3398_/Q sky130_fd_sc_hd__dfxtp_1
X_2418_ hold6/A _2418_/B vssd1 vssd1 vccd1 vccd1 _2507_/C sky130_fd_sc_hd__or2_2
XANTENNA__2874__A1 _2339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2349_ _3377_/Q _2348_/X hold806/X vssd1 vssd1 vccd1 vccd1 _2349_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_47_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2485__S0 _1943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2315__B1_N _2017_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2396__A _2396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1720_ _3533_/Q _1720_/B vssd1 vssd1 vccd1 vccd1 _1720_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 input12/A sky130_fd_sc_hd__dlygate4sd3_1
X_1651_ _3620_/Q hold33/X hold60/X vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__mux2_1
Xhold119 hold119/A vssd1 vssd1 vccd1 vccd1 input27/A sky130_fd_sc_hd__dlygate4sd3_1
X_3321_ _3488_/CLK _3321_/D vssd1 vssd1 vccd1 vccd1 _3321_/Q sky130_fd_sc_hd__dfxtp_1
X_1582_ _1855_/A vssd1 vssd1 vccd1 vccd1 _1582_/Y sky130_fd_sc_hd__inv_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _3331_/CLK _3252_/D vssd1 vssd1 vccd1 vccd1 _3252_/Q sky130_fd_sc_hd__dfxtp_1
X_2203_ _2208_/A _2211_/B vssd1 vssd1 vccd1 vccd1 _2212_/C sky130_fd_sc_hd__nand2_1
X_3183_ _3404_/CLK _3183_/D vssd1 vssd1 vccd1 vccd1 _3183_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2134_ _2134_/A _2134_/B _2134_/C vssd1 vssd1 vccd1 vccd1 _2136_/D sky130_fd_sc_hd__and3_1
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2065_ _2071_/B _2069_/B _2121_/A vssd1 vssd1 vccd1 vccd1 _2068_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_16_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3609_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2967_ _3073_/A vssd1 vssd1 vccd1 vccd1 _2967_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2467__S0 _1943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2792__A0 _2812_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2898_ hold576/X _2101_/X _2904_/S vssd1 vssd1 vccd1 vccd1 _2898_/X sky130_fd_sc_hd__mux2_1
X_1918_ _1911_/B _2554_/S0 _1933_/A vssd1 vssd1 vccd1 vccd1 _1918_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1849_ _1849_/A _1849_/B _1865_/B vssd1 vssd1 vccd1 vccd1 _1850_/A sky130_fd_sc_hd__and3_1
XFILLER_0_71_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold620 _3391_/Q vssd1 vssd1 vccd1 vccd1 hold620/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 _2887_/X vssd1 vssd1 vccd1 vccd1 _3411_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 _3172_/Q vssd1 vssd1 vccd1 vccd1 hold642/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 _2878_/X vssd1 vssd1 vccd1 vccd1 _3403_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 _2614_/X vssd1 vssd1 vccd1 vccd1 _3156_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 _2849_/X vssd1 vssd1 vccd1 vccd1 _3372_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 _3370_/Q vssd1 vssd1 vccd1 vccd1 hold686/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 _3187_/Q vssd1 vssd1 vccd1 vccd1 hold664/X sky130_fd_sc_hd__dlygate4sd3_1
X_3519_ _3623_/CLK _3519_/D _3013_/Y vssd1 vssd1 vccd1 vccd1 _3519_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2783__A0 _2813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3015__A _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2449__S0 _1943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2821_ hold540/X _2075_/B _2823_/S vssd1 vssd1 vccd1 vccd1 _2821_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2752_ _2812_/A1 hold269/X _2753_/S vssd1 vssd1 vccd1 vccd1 _2752_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1703_ _1703_/A _1703_/B vssd1 vssd1 vccd1 vccd1 _1703_/Y sky130_fd_sc_hd__nand2_1
X_2683_ _3492_/Q _3491_/Q _2587_/C vssd1 vssd1 vccd1 vccd1 _2764_/A sky130_fd_sc_hd__or3b_2
X_1634_ _3634_/Q hold2/X hold8/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__mux2_1
X_1565_ _3627_/Q vssd1 vssd1 vccd1 vccd1 _1565_/Y sky130_fd_sc_hd__inv_2
XANTENNA_hold41_A hold41/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3304_ _3488_/CLK _3304_/D vssd1 vssd1 vccd1 vccd1 _3304_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3235_ _3325_/CLK _3235_/D vssd1 vssd1 vccd1 vccd1 _3235_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2829__A1 _2111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3166_ _3433_/CLK _3166_/D vssd1 vssd1 vccd1 vccd1 _3166_/Q sky130_fd_sc_hd__dfxtp_1
X_2117_ hold80/X _2111_/A hold70/X _2115_/A vssd1 vssd1 vccd1 vccd1 _2117_/X sky130_fd_sc_hd__o211a_1
X_3097_ _3105_/A vssd1 vssd1 vccd1 vccd1 _3097_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_55_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2048_ _2047_/X _2046_/X _3489_/Q vssd1 vssd1 vccd1 vccd1 _2049_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout69 _2101_/X vssd1 vssd1 vccd1 vccd1 _2105_/A sky130_fd_sc_hd__buf_4
XANTENNA__2765__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold461 _3295_/Q vssd1 vssd1 vccd1 vccd1 hold461/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 _3484_/Q vssd1 vssd1 vccd1 vccd1 _2205_/A sky130_fd_sc_hd__clkbuf_2
Xhold450 _3214_/Q vssd1 vssd1 vccd1 vccd1 hold450/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 _3519_/Q vssd1 vssd1 vccd1 vccd1 hold483/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _1935_/X vssd1 vssd1 vccd1 vccd1 _3518_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2613__S _2618_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3020_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3020_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2584__A _2585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2804_ _2804_/A _2804_/B vssd1 vssd1 vccd1 vccd1 _2813_/S sky130_fd_sc_hd__nor2_4
XANTENNA__2747__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2735_ _2805_/A1 hold252/X _2743_/S vssd1 vssd1 vccd1 vccd1 _2735_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2666_ _2807_/A1 hold223/X _2672_/S vssd1 vssd1 vccd1 vccd1 _2666_/X sky130_fd_sc_hd__mux2_1
X_1617_ hold28/X hold95/X vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__nand2_2
XFILLER_0_22_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2597_ hold452/X _2813_/A1 _2597_/S vssd1 vssd1 vccd1 vccd1 _2597_/X sky130_fd_sc_hd__mux2_1
X_3218_ _3328_/CLK _3218_/D vssd1 vssd1 vccd1 vccd1 _3218_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_31_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3629_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3149_ _3436_/CLK _3149_/D vssd1 vssd1 vccd1 vccd1 _3149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2433__S _2551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2738__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold280 _3280_/Q vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2910__A0 _2111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold291 _1643_/X vssd1 vssd1 vccd1 vccd1 _3625_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_87_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2729__A0 _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2520_ _2519_/X _2518_/X _3521_/Q vssd1 vssd1 vccd1 vccd1 _2520_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2579__A _2583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2451_ _3369_/Q _3351_/Q _3360_/Q _3189_/Q _2554_/S0 _1911_/B vssd1 vssd1 vccd1 vccd1
+ _2451_/X sky130_fd_sc_hd__mux4_1
X_2382_ hold927/X _2915_/C _1889_/Y vssd1 vssd1 vccd1 vccd1 _2382_/X sky130_fd_sc_hd__a21o_1
Xinput4 input4/A vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_2
X_3003_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3003_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2718_ _2808_/A1 hold154/X _2723_/S vssd1 vssd1 vccd1 vccd1 _2718_/X sky130_fd_sc_hd__mux2_1
X_2649_ _2338_/B hold734/X _2650_/S vssd1 vssd1 vccd1 vccd1 _2649_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2043__S1 _2044_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2399__A hold33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1951_ _2129_/A _3496_/Q vssd1 vssd1 vccd1 vccd1 _1951_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_83_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1882_ _1835_/A _1879_/B _1881_/Y _1838_/B _1560_/Y vssd1 vssd1 vccd1 vccd1 _1882_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3621_ _3629_/CLK _3621_/D _3112_/Y vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__dfrtp_1
X_3552_ _3559_/CLK _3552_/D _3046_/Y vssd1 vssd1 vccd1 vccd1 _3552_/Q sky130_fd_sc_hd__dfrtp_1
X_2503_ _3183_/Q _3336_/Q _3165_/Q _3147_/Q _1943_/B _2550_/S1 vssd1 vssd1 vccd1 vccd1
+ _2503_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_3_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3483_ _3483_/CLK _3483_/D _2977_/Y vssd1 vssd1 vccd1 vccd1 _3483_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2025__S1 _2222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2434_ _2433_/X _2430_/X _3522_/Q vssd1 vssd1 vccd1 vccd1 _2434_/X sky130_fd_sc_hd__mux2_1
X_2365_ _2365_/A _2365_/B vssd1 vssd1 vccd1 vccd1 _2365_/Y sky130_fd_sc_hd__nor2_1
X_2296_ hold46/X hold41/X hold30/X vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__mux2_1
XANTENNA__1660__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2711__S _2713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1916__A1 _2551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1997__S _2052_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap77 _2597_/S vssd1 vssd1 vccd1 vccd1 _2594_/S sky130_fd_sc_hd__buf_4
XFILLER_0_57_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2621__S _2629_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3018__A _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2150_ _1956_/B _2149_/X _2375_/A vssd1 vssd1 vccd1 vccd1 _2150_/X sky130_fd_sc_hd__o21a_1
X_2081_ _2054_/A _2081_/B _2081_/C vssd1 vssd1 vccd1 vccd1 _2081_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_88_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2983_ _3126_/A vssd1 vssd1 vccd1 vccd1 _2983_/Y sky130_fd_sc_hd__inv_2
X_1934_ _1929_/A _1930_/X _1931_/X _1933_/Y vssd1 vssd1 vccd1 vccd1 _1934_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_83_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1865_ _1865_/A _1865_/B vssd1 vssd1 vccd1 vccd1 _1865_/X sky130_fd_sc_hd__or2_1
Xhold802 _3155_/Q vssd1 vssd1 vccd1 vccd1 hold802/X sky130_fd_sc_hd__dlygate4sd3_1
X_1796_ _1604_/Y _2383_/C _1775_/B _1795_/Y _1794_/X vssd1 vssd1 vccd1 vccd1 _1803_/B
+ sky130_fd_sc_hd__o221a_2
X_3604_ _3604_/CLK _3604_/D _3095_/Y vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__dfrtp_1
X_3535_ _3539_/CLK _3535_/D _3029_/Y vssd1 vssd1 vccd1 vccd1 _3535_/Q sky130_fd_sc_hd__dfrtp_1
Xhold846 _1882_/X vssd1 vssd1 vccd1 vccd1 _3529_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 _2234_/Y vssd1 vssd1 vccd1 vccd1 _3481_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold813 _2252_/X vssd1 vssd1 vccd1 vccd1 _3474_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold824 _3509_/Q vssd1 vssd1 vccd1 vccd1 hold824/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold868 _1880_/X vssd1 vssd1 vccd1 vccd1 _3530_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 _3584_/Q vssd1 vssd1 vccd1 vccd1 hold857/X sky130_fd_sc_hd__dlygate4sd3_1
X_3466_ _3579_/CLK _3466_/D _2960_/Y vssd1 vssd1 vccd1 vccd1 _3466_/Q sky130_fd_sc_hd__dfrtp_4
Xhold879 _3559_/Q vssd1 vssd1 vccd1 vccd1 _1778_/A sky130_fd_sc_hd__buf_1
X_2417_ _3594_/Q _2417_/B vssd1 vssd1 vccd1 vccd1 _2417_/X sky130_fd_sc_hd__or2_1
XFILLER_0_58_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3397_ _3433_/CLK _3397_/D vssd1 vssd1 vccd1 vccd1 _3397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2348_ _1570_/Y _2105_/B _2344_/X _2345_/X _2347_/Y vssd1 vssd1 vccd1 vccd1 _2348_/X
+ sky130_fd_sc_hd__o2111a_1
X_2279_ _3462_/Q _2283_/B _2273_/A vssd1 vssd1 vccd1 vccd1 _2279_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__2706__S _2713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2485__S1 _2550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2562__A1 _2506_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2616__S _2618_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuart_macro_wrapper_131 vssd1 vssd1 vccd1 vccd1 uart_macro_wrapper_131/HI io_oeb[1]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1650_ hold87/X hold52/X hold60/X vssd1 vssd1 vccd1 vccd1 _3621_/D sky130_fd_sc_hd__mux2_1
X_1581_ _3543_/Q vssd1 vssd1 vccd1 vccd1 _1581_/Y sky130_fd_sc_hd__inv_2
Xhold109 _1624_/C vssd1 vssd1 vccd1 vccd1 _1657_/C sky130_fd_sc_hd__dlygate4sd3_1
X_3320_ _3488_/CLK _3320_/D vssd1 vssd1 vccd1 vccd1 _3320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2305__A1 _2396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3330_/CLK _3251_/D vssd1 vssd1 vccd1 vccd1 _3251_/Q sky130_fd_sc_hd__dfxtp_1
X_3182_ _3404_/CLK _3182_/D vssd1 vssd1 vccd1 vccd1 _3182_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2202_ _2202_/A _2202_/B vssd1 vssd1 vccd1 vccd1 _2214_/B sky130_fd_sc_hd__nand2_2
X_2133_ _2366_/A _2133_/B _2133_/C _2133_/D vssd1 vssd1 vccd1 vccd1 _2136_/C sky130_fd_sc_hd__and4_2
X_2064_ _3550_/Q _2089_/B vssd1 vssd1 vccd1 vccd1 _2069_/B sky130_fd_sc_hd__nand2_1
X_2966_ _3073_/A vssd1 vssd1 vccd1 vccd1 _2966_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2467__S1 _2550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2897_ hold570/X _2091_/X _2904_/S vssd1 vssd1 vccd1 vccd1 _2897_/X sky130_fd_sc_hd__mux2_1
X_1917_ _1933_/A _1909_/B _1911_/C vssd1 vssd1 vccd1 vccd1 _1917_/X sky130_fd_sc_hd__o21a_1
X_1848_ _1865_/A _1865_/B vssd1 vssd1 vccd1 vccd1 _1848_/Y sky130_fd_sc_hd__nand2_1
Xhold610 _3160_/Q vssd1 vssd1 vccd1 vccd1 hold610/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 _2864_/X vssd1 vssd1 vccd1 vccd1 _3391_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 _3180_/Q vssd1 vssd1 vccd1 vccd1 hold654/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold632 _3162_/Q vssd1 vssd1 vccd1 vccd1 hold632/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 _2634_/X vssd1 vssd1 vccd1 vccd1 _3172_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1779_ _3625_/Q _3624_/Q vssd1 vssd1 vccd1 vccd1 _1784_/A sky130_fd_sc_hd__nor2_1
Xhold687 _2847_/X vssd1 vssd1 vccd1 vccd1 _3370_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 _3152_/Q vssd1 vssd1 vccd1 vccd1 hold676/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 _2650_/X vssd1 vssd1 vccd1 vccd1 _3187_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3518_ _3623_/CLK _3518_/D _3012_/Y vssd1 vssd1 vccd1 vccd1 _3518_/Q sky130_fd_sc_hd__dfrtp_1
X_3449_ _3633_/CLK hold73/X _2943_/Y vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__dfrtp_1
Xhold698 _3362_/Q vssd1 vssd1 vccd1 vccd1 hold698/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1969__S0 _2224_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2535__A1 _2583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2535__B2 _2506_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2820_ hold622/X _2079_/A _2823_/S vssd1 vssd1 vccd1 vccd1 _2820_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2449__S1 _2550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2751_ _2811_/A1 hold368/X _2753_/S vssd1 vssd1 vccd1 vccd1 _2751_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1702_ _1700_/C hold898/X _3466_/D vssd1 vssd1 vccd1 vccd1 _1702_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2682_ hold450/X _2813_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2682_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_81_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1633_ _3635_/Q hold41/X hold8/X vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1564_ hold90/X vssd1 vssd1 vccd1 vccd1 _2115_/A sky130_fd_sc_hd__inv_2
X_3303_ _3488_/CLK _3303_/D vssd1 vssd1 vccd1 vccd1 _3303_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2110__A _2111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3234_ _3328_/CLK _3234_/D vssd1 vssd1 vccd1 vccd1 _3234_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3165_ _3404_/CLK _3165_/D vssd1 vssd1 vccd1 vccd1 _3165_/Q sky130_fd_sc_hd__dfxtp_1
X_3096_ _3124_/A vssd1 vssd1 vccd1 vccd1 _3096_/Y sky130_fd_sc_hd__inv_2
X_2116_ hold70/X _2116_/B _2115_/Y vssd1 vssd1 vccd1 vccd1 _2116_/X sky130_fd_sc_hd__or3b_1
X_2047_ _3242_/Q _3314_/Q _3305_/Q _3296_/Q _1590_/A _2222_/A vssd1 vssd1 vccd1 vccd1
+ _2047_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2949_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2949_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold462 _2773_/X vssd1 vssd1 vccd1 vccd1 _3295_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 _2682_/X vssd1 vssd1 vccd1 vccd1 _3214_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold440 _3232_/Q vssd1 vssd1 vccd1 vccd1 hold440/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 _2219_/X vssd1 vssd1 vccd1 vccd1 _3484_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 _1920_/X vssd1 vssd1 vccd1 vccd1 _3519_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 hold495/A vssd1 vssd1 vccd1 vccd1 _2145_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_67_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2756__A1 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_1_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3436_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2692__A0 _2812_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2803_ hold463/X _2813_/A1 _2803_/S vssd1 vssd1 vccd1 vccd1 _2803_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2105__A _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2734_ _2804_/A _2794_/A _2794_/B vssd1 vssd1 vccd1 vccd1 _2743_/S sky130_fd_sc_hd__or3b_4
X_2665_ _2806_/A1 hold159/X _2672_/S vssd1 vssd1 vccd1 vccd1 _2665_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2596_ hold345/X _2812_/A1 _2597_/S vssd1 vssd1 vccd1 vccd1 _2596_/X sky130_fd_sc_hd__mux2_1
X_1616_ hold28/A hold95/A vssd1 vssd1 vccd1 vccd1 _2511_/A sky130_fd_sc_hd__and2_2
X_3217_ _3325_/CLK _3217_/D vssd1 vssd1 vccd1 vccd1 _3217_/Q sky130_fd_sc_hd__dfxtp_1
X_3148_ _3433_/CLK _3148_/D vssd1 vssd1 vccd1 vccd1 _3148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3079_ _3133_/A vssd1 vssd1 vccd1 vccd1 _3079_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_72_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold492_A _3522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold270 _2752_/X vssd1 vssd1 vccd1 vccd1 _3276_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold281 _2757_/X vssd1 vssd1 vccd1 vccd1 _3280_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _3294_/Q vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2624__S _2629_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2450_ _2449_/X _2448_/X _2551_/S vssd1 vssd1 vccd1 vccd1 _2450_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2381_ _2381_/A _2381_/B vssd1 vssd1 vccd1 vccd1 _2915_/C sky130_fd_sc_hd__nand2_1
Xinput5 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_1
XANTENNA__2665__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3002_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3002_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_36_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2534__S _3522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1640__A1 hold86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout126_A _3131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2717_ _2807_/A1 hold217/X _2723_/S vssd1 vssd1 vccd1 vccd1 _2717_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2648_ _2075_/B hold772/X _2650_/S vssd1 vssd1 vccd1 vccd1 _2648_/X sky130_fd_sc_hd__mux2_1
X_2579_ _2583_/B _2579_/B vssd1 vssd1 vccd1 vccd1 _2579_/X sky130_fd_sc_hd__and2_1
XFILLER_0_10_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2709__S _2713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2656__A0 _2111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2503__S0 _1943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2647__A0 _2079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1950_ _2367_/A _1950_/B vssd1 vssd1 vccd1 vccd1 _2366_/A sky130_fd_sc_hd__nor2_2
X_1881_ _1881_/A _1881_/B vssd1 vssd1 vccd1 vccd1 _1881_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__1622__A1 _2395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3620_ _3623_/CLK hold61/X _3111_/Y vssd1 vssd1 vccd1 vccd1 _3620_/Q sky130_fd_sc_hd__dfrtp_1
X_3551_ _3551_/CLK _3551_/D _3045_/Y vssd1 vssd1 vccd1 vccd1 _3551_/Q sky130_fd_sc_hd__dfrtp_1
X_2502_ _3405_/Q _3396_/Q _3387_/Q _3432_/Q _1943_/B _2550_/S1 vssd1 vssd1 vccd1 vccd1
+ _2502_/X sky130_fd_sc_hd__mux4_1
X_3482_ _3610_/CLK _3482_/D _2976_/Y vssd1 vssd1 vccd1 vccd1 _3482_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2433_ _2432_/X _2431_/X _2551_/S vssd1 vssd1 vccd1 vccd1 _2433_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1689__A1 _2395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2364_ _2361_/X _2362_/X _2363_/X _1598_/Y vssd1 vssd1 vccd1 vccd1 _2365_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2295_ _3456_/Q hold76/X hold30/X vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__mux2_1
XANTENNA__1660__C input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2638__A0 _2075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2877__A0 _2097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2341__A2 _2079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2629__A0 _2339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2902__S _2904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2332__A2 _1889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2080_ _2080_/A _2080_/B vssd1 vssd1 vccd1 vccd1 _2081_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2982_ _3126_/A vssd1 vssd1 vccd1 vccd1 _2982_/Y sky130_fd_sc_hd__inv_2
X_1933_ _1933_/A _1933_/B vssd1 vssd1 vccd1 vccd1 _1933_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2812__S _2813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1864_ _1835_/A _1851_/B _1863_/X _1849_/A _1560_/Y vssd1 vssd1 vccd1 vccd1 _1864_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_71_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput30 hold85/X vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__clkbuf_2
X_3603_ _3604_/CLK _3603_/D _3094_/Y vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__dfrtp_1
Xhold803 _2613_/X vssd1 vssd1 vccd1 vccd1 _3155_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1795_ _1815_/B _1795_/B vssd1 vssd1 vccd1 vccd1 _1795_/Y sky130_fd_sc_hd__nand2_1
X_3534_ _3539_/CLK _3534_/D _3028_/Y vssd1 vssd1 vccd1 vccd1 _3534_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold836 _3546_/Q vssd1 vssd1 vccd1 vccd1 hold836/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 _3508_/Q vssd1 vssd1 vccd1 vccd1 hold814/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 _2009_/X vssd1 vssd1 vccd1 vccd1 _3509_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3465_ _3637_/CLK _3465_/D _2959_/Y vssd1 vssd1 vccd1 vccd1 _3465_/Q sky130_fd_sc_hd__dfrtp_1
Xhold847 _3593_/Q vssd1 vssd1 vccd1 vccd1 hold847/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 _1691_/X vssd1 vssd1 vccd1 vccd1 _3594_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 _3585_/Q vssd1 vssd1 vccd1 vccd1 hold869/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2859__A0 _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2416_ _2416_/A _2568_/C vssd1 vssd1 vccd1 vccd1 _2417_/B sky130_fd_sc_hd__and2_2
X_3396_ _3435_/CLK _3396_/D vssd1 vssd1 vccd1 vccd1 _3396_/Q sky130_fd_sc_hd__dfxtp_1
X_2347_ hold288/X _2092_/Y _2110_/Y hold105/X _2346_/X vssd1 vssd1 vccd1 vccd1 _2347_/Y
+ sky130_fd_sc_hd__a221oi_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2278_ _2285_/A _2278_/B _2278_/C vssd1 vssd1 vccd1 vccd1 _2278_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_74_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2632__S _2640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuart_macro_wrapper_132 vssd1 vssd1 vccd1 vccd1 uart_macro_wrapper_132/HI wbs_dat_o[17]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1580_ _1580_/A vssd1 vssd1 vccd1 vccd1 _1817_/A sky130_fd_sc_hd__inv_2
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3483_/CLK _3250_/D vssd1 vssd1 vccd1 vccd1 _3250_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _3414_/CLK _3181_/D vssd1 vssd1 vccd1 vccd1 _3181_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _2214_/A _2201_/B _2211_/B vssd1 vssd1 vccd1 vccd1 _2202_/B sky130_fd_sc_hd__or3b_1
X_2132_ _2149_/A _2366_/B _3346_/Q vssd1 vssd1 vccd1 vccd1 _2133_/D sky130_fd_sc_hd__mux2_1
XANTENNA__2807__S _2813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2063_ _3551_/Q _2089_/B vssd1 vssd1 vccd1 vccd1 _2071_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_76_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2965_ _3073_/A vssd1 vssd1 vccd1 vccd1 _2965_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2896_ hold612/X _2096_/Y _2904_/S vssd1 vssd1 vccd1 vccd1 _2896_/X sky130_fd_sc_hd__mux2_1
X_1916_ _2551_/S _1910_/B _1910_/Y _2164_/B vssd1 vssd1 vccd1 vccd1 _3521_/D sky130_fd_sc_hd__a22o_1
X_1847_ _1847_/A _1847_/B vssd1 vssd1 vccd1 vccd1 _1865_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_25_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3542_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold600 _3173_/Q vssd1 vssd1 vccd1 vccd1 hold600/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold611 _2618_/X vssd1 vssd1 vccd1 vccd1 _3160_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold622 _3337_/Q vssd1 vssd1 vccd1 vccd1 hold622/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 _3195_/Q vssd1 vssd1 vccd1 vccd1 hold644/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 _2622_/X vssd1 vssd1 vccd1 vccd1 _3162_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1778_ _1778_/A _2321_/B vssd1 vssd1 vccd1 vccd1 _1792_/B sky130_fd_sc_hd__xnor2_1
X_3517_ _3623_/CLK _3517_/D _3011_/Y vssd1 vssd1 vccd1 vccd1 _3517_/Q sky130_fd_sc_hd__dfrtp_1
Xhold677 _2610_/X vssd1 vssd1 vccd1 vccd1 _3152_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 _3369_/Q vssd1 vssd1 vccd1 vccd1 hold688/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 _2643_/X vssd1 vssd1 vccd1 vccd1 _3180_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 _3167_/Q vssd1 vssd1 vccd1 vccd1 hold666/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 _2838_/X vssd1 vssd1 vccd1 vccd1 _3362_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3448_ _3642_/CLK hold89/X _2942_/Y vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__dfrtp_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ _3642_/CLK _3379_/D _2927_/Y vssd1 vssd1 vccd1 vccd1 _3379_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_3__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__1969__S1 _2193_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2299__A1 hold49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2200__B _2200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2627__S _2629_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2750_ _2810_/A1 hold331/X _2753_/S vssd1 vssd1 vccd1 vccd1 _2750_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1701_ _1701_/A _1701_/B vssd1 vssd1 vccd1 vccd1 _1701_/Y sky130_fd_sc_hd__nand2_1
X_2681_ hold376/X _2812_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2681_/X sky130_fd_sc_hd__mux2_1
X_1632_ _2263_/A hold76/X hold8/X vssd1 vssd1 vccd1 vccd1 _1632_/X sky130_fd_sc_hd__mux2_1
X_1563_ hold54/X vssd1 vssd1 vccd1 vccd1 _1563_/Y sky130_fd_sc_hd__inv_2
X_3302_ _3488_/CLK _3302_/D vssd1 vssd1 vccd1 vccd1 _3302_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _3330_/CLK _3233_/D vssd1 vssd1 vccd1 vccd1 _3233_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3164_ _3404_/CLK _3164_/D vssd1 vssd1 vccd1 vccd1 _3164_/Q sky130_fd_sc_hd__dfxtp_1
X_3095_ _3095_/A vssd1 vssd1 vccd1 vccd1 _3095_/Y sky130_fd_sc_hd__inv_2
X_2115_ _2115_/A hold80/X vssd1 vssd1 vccd1 vccd1 _2115_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_55_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2046_ _3287_/Q _3278_/Q _3269_/Q _3260_/Q _1590_/A _2222_/A vssd1 vssd1 vccd1 vccd1
+ _2046_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_9_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1677__A hold65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2948_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2948_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_72_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2879_ _2105_/B hold722/X _2884_/S vssd1 vssd1 vccd1 vccd1 _2879_/X sky130_fd_sc_hd__mux2_1
Xhold463 _3322_/Q vssd1 vssd1 vccd1 vccd1 hold463/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 _3142_/Q vssd1 vssd1 vccd1 vccd1 hold452/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold430 _3139_/Q vssd1 vssd1 vccd1 vccd1 hold430/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 _2703_/X vssd1 vssd1 vccd1 vccd1 _3232_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 _3485_/Q vssd1 vssd1 vccd1 vccd1 _2208_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold485 _3495_/Q vssd1 vssd1 vccd1 vccd1 _1921_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 _2200_/B vssd1 vssd1 vccd1 vccd1 _2375_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2910__S _2914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2141__B1 _2052_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2802_ hold294/X _2812_/A1 _2803_/S vssd1 vssd1 vccd1 vccd1 _2802_/X sky130_fd_sc_hd__mux2_1
X_2733_ _2813_/A1 hold442/X _2733_/S vssd1 vssd1 vccd1 vccd1 _2733_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2105__B _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2664_ _2805_/A1 hold239/X _2672_/S vssd1 vssd1 vccd1 vccd1 _2664_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2595_ hold445/X _2811_/A1 _2597_/S vssd1 vssd1 vccd1 vccd1 _2595_/X sky130_fd_sc_hd__mux2_1
X_1615_ hold18/X hold58/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__nor2_1
XFILLER_0_5_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3216_ _3331_/CLK _3216_/D vssd1 vssd1 vccd1 vccd1 _3216_/Q sky130_fd_sc_hd__dfxtp_1
X_3147_ _3404_/CLK _3147_/D vssd1 vssd1 vccd1 vccd1 _3147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3078_ _3105_/A vssd1 vssd1 vccd1 vccd1 _3078_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_82_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2029_ _2029_/A vssd1 vssd1 vccd1 vccd1 _2029_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2435__A1 _2506_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3416_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1946__B1 _2551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2046__S0 _1590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold271 _3611_/Q vssd1 vssd1 vccd1 vccd1 _1575_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold260 _2177_/X vssd1 vssd1 vccd1 vccd1 _3493_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 _2772_/X vssd1 vssd1 vccd1 vccd1 _3294_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _3224_/Q vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2674__A1 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2640__S _2640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2380_ _2187_/A _1956_/B _2367_/X _2149_/A vssd1 vssd1 vccd1 vccd1 _3347_/D sky130_fd_sc_hd__a22o_1
Xinput6 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
X_3001_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3001_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1955__A _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2716_ _2806_/A1 hold171/X _2723_/S vssd1 vssd1 vccd1 vccd1 _2716_/X sky130_fd_sc_hd__mux2_1
X_2647_ _2079_/A hold792/X _2650_/S vssd1 vssd1 vccd1 vccd1 _2647_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2578_ _2511_/Y _2581_/C _2577_/X _2511_/B _3457_/Q vssd1 vssd1 vccd1 vccd1 _2579_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2503__S1 _2550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2635__S _2640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1880_ _1835_/A _1839_/Y _1879_/Y _1838_/A _1560_/Y vssd1 vssd1 vccd1 vccd1 _1880_/X
+ sky130_fd_sc_hd__a32o_1
X_3550_ _3551_/CLK _3550_/D _3044_/Y vssd1 vssd1 vccd1 vccd1 _3550_/Q sky130_fd_sc_hd__dfrtp_1
X_2501_ _2500_/X _2499_/X _3521_/Q vssd1 vssd1 vccd1 vccd1 _2501_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3481_ _3499_/CLK _3481_/D _2975_/Y vssd1 vssd1 vccd1 vccd1 _3481_/Q sky130_fd_sc_hd__dfrtp_1
X_2432_ _3170_/Q _3419_/Q _3410_/Q _3152_/Q _1911_/C _1911_/B vssd1 vssd1 vccd1 vccd1
+ _2432_/X sky130_fd_sc_hd__mux4_1
X_2363_ _3571_/Q _3570_/Q _3569_/Q _3568_/Q vssd1 vssd1 vccd1 vccd1 _2363_/X sky130_fd_sc_hd__or4_1
X_2294_ _3457_/Q hold36/X hold30/X vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__mux2_1
XANTENNA__1660__D input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2810__A1 _2810_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap79 _2381_/A vssd1 vssd1 vccd1 vccd1 _1795_/B sky130_fd_sc_hd__buf_2
XANTENNA__2488__S0 _2554_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2801__A1 _2811_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2868__A1 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2981_ _3126_/A vssd1 vssd1 vccd1 vccd1 _2981_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1932_ _1929_/A _1930_/X _1931_/X vssd1 vssd1 vccd1 vccd1 _1932_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1863_ _3537_/Q _3536_/Q _1846_/A _1849_/A vssd1 vssd1 vccd1 vccd1 _1863_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3602_ _3633_/CLK _3602_/D _3093_/Y vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__dfrtp_1
Xinput31 hold32/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__buf_1
Xinput20 input20/A vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1794_ _1815_/B _1795_/B _1794_/A3 _1793_/Y _1824_/A vssd1 vssd1 vccd1 vccd1 _1794_/X
+ sky130_fd_sc_hd__a32o_1
X_3533_ _3539_/CLK _3533_/D _3027_/Y vssd1 vssd1 vccd1 vccd1 _3533_/Q sky130_fd_sc_hd__dfrtp_1
Xhold826 _3583_/Q vssd1 vssd1 vccd1 vccd1 hold826/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 _1831_/X vssd1 vssd1 vccd1 vccd1 _3545_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold804 _3383_/Q vssd1 vssd1 vccd1 vccd1 hold804/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold57_A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold815 _2020_/X vssd1 vssd1 vccd1 vccd1 _3508_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3464_ _3637_/CLK _3464_/D _2958_/Y vssd1 vssd1 vccd1 vccd1 _3464_/Q sky130_fd_sc_hd__dfrtp_1
Xhold848 _2331_/X vssd1 vssd1 vccd1 vccd1 _3381_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold859 _3547_/Q vssd1 vssd1 vccd1 vccd1 hold859/X sky130_fd_sc_hd__dlygate4sd3_1
X_2415_ _2415_/A _2419_/B vssd1 vssd1 vccd1 vccd1 _2568_/C sky130_fd_sc_hd__nand2_2
X_3395_ _3433_/CLK _3395_/D vssd1 vssd1 vccd1 vccd1 _3395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2346_ hold288/X _2092_/Y _2105_/A _1571_/Y vssd1 vssd1 vccd1 vccd1 _2346_/X sky130_fd_sc_hd__a2bb2o_1
X_2277_ _2277_/A _2280_/B vssd1 vssd1 vccd1 vccd1 _2278_/C sky130_fd_sc_hd__or2_1
XFILLER_0_74_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_2__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_2__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__1770__A1 _3443_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2913__S _2914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2786__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xuart_macro_wrapper_133 vssd1 vssd1 vccd1 vccd1 uart_macro_wrapper_133/HI wbs_dat_o[20]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_80_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _2661_/B _2200_/B vssd1 vssd1 vccd1 vccd1 _2211_/B sky130_fd_sc_hd__nand2_2
X_3180_ _3414_/CLK _3180_/D vssd1 vssd1 vccd1 vccd1 _3180_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2710__A0 _2810_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2131_ _2149_/A _2367_/C vssd1 vssd1 vccd1 vccd1 _2133_/C sky130_fd_sc_hd__nand2_1
X_2062_ _2071_/A _2062_/B vssd1 vssd1 vccd1 vccd1 _2062_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2964_ _3073_/A vssd1 vssd1 vccd1 vccd1 _2964_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2777__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1915_ _1915_/A _1915_/B vssd1 vssd1 vccd1 vccd1 _2164_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_29_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2895_ _3526_/Q _2905_/B _2895_/C vssd1 vssd1 vccd1 vccd1 _2904_/S sky130_fd_sc_hd__nor3_4
X_1846_ _1846_/A vssd1 vssd1 vccd1 vccd1 _1847_/B sky130_fd_sc_hd__inv_2
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold601 _2635_/X vssd1 vssd1 vccd1 vccd1 _3173_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold612 _3419_/Q vssd1 vssd1 vccd1 vccd1 hold612/X sky130_fd_sc_hd__dlygate4sd3_1
X_1777_ _2121_/A _2056_/A _3627_/Q vssd1 vssd1 vccd1 vccd1 _2321_/B sky130_fd_sc_hd__o21a_1
Xhold623 _2820_/X vssd1 vssd1 vccd1 vccd1 _3337_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 _2659_/X vssd1 vssd1 vccd1 vccd1 _3195_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 _3376_/Q vssd1 vssd1 vccd1 vccd1 hold634/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout101_A hold49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3516_ _3612_/CLK _3516_/D _3010_/Y vssd1 vssd1 vccd1 vccd1 _3516_/Q sky130_fd_sc_hd__dfrtp_1
Xhold667 _2627_/X vssd1 vssd1 vccd1 vccd1 _3167_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold678 _3169_/Q vssd1 vssd1 vccd1 vccd1 hold678/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 _3425_/Q vssd1 vssd1 vccd1 vccd1 hold656/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold689 _2846_/X vssd1 vssd1 vccd1 vccd1 _3369_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3447_ _3642_/CLK _3447_/D _2941_/Y vssd1 vssd1 vccd1 vccd1 _3447_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ _3633_/CLK _3378_/D _2926_/Y vssd1 vssd1 vccd1 vccd1 _3378_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2701__A0 _2811_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2329_ _2145_/D _2326_/X hold891/X vssd1 vssd1 vccd1 vccd1 _3443_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_39_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2465__C1 _2583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2018__B _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2768__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2908__S _2914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1700_ _1700_/A _1700_/B _1700_/C vssd1 vssd1 vccd1 vccd1 _1700_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_30_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2680_ hold432/X _2811_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2680_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1631_ hold38/X hold36/X hold8/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__mux2_1
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1562_ _3634_/Q vssd1 vssd1 vccd1 vccd1 _2567_/A sky130_fd_sc_hd__inv_2
X_3301_ _3305_/CLK _3301_/D vssd1 vssd1 vccd1 vccd1 _3301_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ _3513_/CLK _3232_/D vssd1 vssd1 vccd1 vccd1 _3232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ _3414_/CLK _3163_/D vssd1 vssd1 vccd1 vccd1 _3163_/Q sky130_fd_sc_hd__dfxtp_1
X_2114_ hold70/X _2116_/B _2114_/C vssd1 vssd1 vccd1 vccd1 _2114_/Y sky130_fd_sc_hd__nand3b_1
X_3094_ _3095_/A vssd1 vssd1 vccd1 vccd1 _3094_/Y sky130_fd_sc_hd__inv_2
X_2045_ _2043_/X _2044_/X _2045_/S vssd1 vssd1 vccd1 vccd1 _2045_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2447__C1 _2583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2947_ _3128_/A vssd1 vssd1 vccd1 vccd1 _2947_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2878_ _2105_/A hold630/X _2884_/S vssd1 vssd1 vccd1 vccd1 _2878_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1829_ hold861/X hold859/X _1831_/S vssd1 vssd1 vccd1 vccd1 _1829_/X sky130_fd_sc_hd__mux2_1
Xhold420 _3246_/Q vssd1 vssd1 vccd1 vccd1 hold420/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 _3259_/Q vssd1 vssd1 vccd1 vccd1 hold442/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 _2597_/X vssd1 vssd1 vccd1 vccd1 _3142_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold431 _2594_/X vssd1 vssd1 vccd1 vccd1 _3139_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 _2803_/X vssd1 vssd1 vccd1 vccd1 _3322_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 _2217_/X vssd1 vssd1 vccd1 vccd1 _3485_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 _1919_/X vssd1 vssd1 vccd1 vccd1 _3520_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold497 _2188_/Y vssd1 vssd1 vccd1 vccd1 _2196_/B sky130_fd_sc_hd__buf_1
XANTENNA__1632__S hold8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2913__A0 _2338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2638__S _2640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2801_ hold386/X _2811_/A1 _2803_/S vssd1 vssd1 vccd1 vccd1 _2801_/X sky130_fd_sc_hd__mux2_1
X_2732_ _2812_/A1 hold408/X _2733_/S vssd1 vssd1 vccd1 vccd1 _2732_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2663_ _2784_/C _2804_/B vssd1 vssd1 vccd1 vccd1 _2672_/S sky130_fd_sc_hd__or2_4
X_2594_ hold430/X _2810_/A1 _2594_/S vssd1 vssd1 vccd1 vccd1 _2594_/X sky130_fd_sc_hd__mux2_1
X_1614_ _2287_/A hold57/X _1624_/C hold5/X vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__or4bb_1
XANTENNA__2402__A hold49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3215_ _3325_/CLK _3215_/D vssd1 vssd1 vccd1 vccd1 _3215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3146_ _3404_/CLK _3146_/D vssd1 vssd1 vccd1 vccd1 _3146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3077_ _3126_/A vssd1 vssd1 vccd1 vccd1 _3077_/Y sky130_fd_sc_hd__inv_2
X_2028_ _1985_/S _2023_/X _2027_/X vssd1 vssd1 vccd1 vccd1 _2029_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1907__D_N _2506_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold109_A _1624_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2046__S1 _2222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold250 _3298_/Q vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 _3206_/Q vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 _3321_/Q vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2371__A1 _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold272 _3253_/Q vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 _2695_/X vssd1 vssd1 vccd1 vccd1 _3224_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2982__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1598__A _3341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2222__A _2222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 input7/A vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
X_3000_ _3114_/A vssd1 vssd1 vccd1 vccd1 _3000_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2715_ _2805_/A1 hold225/X _2723_/S vssd1 vssd1 vccd1 vccd1 _2715_/X sky130_fd_sc_hd__mux2_1
X_2646_ _2111_/B hold640/X _2650_/S vssd1 vssd1 vccd1 vccd1 _2646_/X sky130_fd_sc_hd__mux2_1
X_2577_ hold38/A hold7/A vssd1 vssd1 vccd1 vccd1 _2577_/X sky130_fd_sc_hd__or2_1
X_3129_ _3133_/A vssd1 vssd1 vccd1 vccd1 _3129_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1919__A1 _1911_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2592__A1 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2977__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3480_ _3571_/CLK _3480_/D _2974_/Y vssd1 vssd1 vccd1 vccd1 _3480_/Q sky130_fd_sc_hd__dfrtp_1
X_2500_ _3174_/Q _3423_/Q _3414_/Q _3156_/Q _2554_/S0 _1911_/B vssd1 vssd1 vccd1 vccd1
+ _2500_/X sky130_fd_sc_hd__mux4_1
X_2431_ _3368_/Q _3350_/Q _3359_/Q _3188_/Q _1911_/C _1942_/A vssd1 vssd1 vccd1 vccd1
+ _2431_/X sky130_fd_sc_hd__mux4_1
X_2362_ _3567_/Q _3566_/Q _3565_/Q _3564_/Q vssd1 vssd1 vccd1 vccd1 _2362_/X sky130_fd_sc_hd__or4_1
X_2293_ _3458_/Q hold11/X hold30/A vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__mux2_1
XFILLER_0_2_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_1__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_19_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3604_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1966__A _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2629_ _2339_/B hold678/X _2629_/S vssd1 vssd1 vccd1 vccd1 _2629_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1640__S hold8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2488__S1 _1911_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1999__S0 _2044_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2317__A1 _2029_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2049__A_N _1985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2980_ _3126_/A vssd1 vssd1 vccd1 vccd1 _2980_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_33_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1931_ _1931_/A _1931_/B vssd1 vssd1 vccd1 vccd1 _1931_/X sky130_fd_sc_hd__xor2_1
X_1862_ _1861_/Y _1859_/B _1583_/A _1560_/Y vssd1 vssd1 vccd1 vccd1 _1862_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_71_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput21 hold1/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__clkbuf_1
Xinput10 input10/A vssd1 vssd1 vccd1 vccd1 _2287_/A sky130_fd_sc_hd__clkbuf_2
X_3601_ _3604_/CLK _3601_/D _3092_/Y vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__dfrtp_1
Xinput32 hold51/X vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__buf_1
X_1793_ _1793_/A vssd1 vssd1 vccd1 vccd1 _1793_/Y sky130_fd_sc_hd__inv_2
X_3532_ _3539_/CLK _3532_/D _3026_/Y vssd1 vssd1 vccd1 vccd1 _3532_/Q sky130_fd_sc_hd__dfrtp_1
Xhold827 _2259_/X vssd1 vssd1 vccd1 vccd1 _3467_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold805 _2856_/X vssd1 vssd1 vccd1 vccd1 _3383_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold816 _3510_/Q vssd1 vssd1 vccd1 vccd1 hold816/X sky130_fd_sc_hd__dlygate4sd3_1
X_3463_ _3637_/CLK _3463_/D _2957_/Y vssd1 vssd1 vccd1 vccd1 _3463_/Q sky130_fd_sc_hd__dfrtp_1
Xhold838 _3579_/Q vssd1 vssd1 vccd1 vccd1 _1700_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 _3478_/Q vssd1 vssd1 vccd1 vccd1 _2260_/B sky130_fd_sc_hd__dlygate4sd3_1
X_2414_ _3584_/Q hold67/A vssd1 vssd1 vccd1 vccd1 _2414_/X sky130_fd_sc_hd__or2_1
X_3394_ _3403_/CLK _3394_/D vssd1 vssd1 vccd1 vccd1 _3394_/Q sky130_fd_sc_hd__dfxtp_1
X_2345_ _1570_/Y _2105_/B _2110_/Y hold105/X vssd1 vssd1 vccd1 vccd1 _2345_/X sky130_fd_sc_hd__o2bb2a_1
X_2276_ _2285_/A _2276_/B vssd1 vssd1 vccd1 vccd1 _2276_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2795__A1 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1635__S hold8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2483__B1 _2583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuart_macro_wrapper_134 vssd1 vssd1 vccd1 vccd1 uart_macro_wrapper_134/HI wbs_dat_o[22]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2130_ _2130_/A _2130_/B _2130_/C vssd1 vssd1 vccd1 vccd1 _2367_/C sky130_fd_sc_hd__or3_1
X_2061_ _3548_/Q _2089_/B vssd1 vssd1 vccd1 vccd1 _2062_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_44_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2963_ _3073_/A vssd1 vssd1 vccd1 vccd1 _2963_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1914_ _1911_/B _1911_/C _1911_/A vssd1 vssd1 vccd1 vccd1 _1915_/B sky130_fd_sc_hd__a21oi_1
X_2894_ _2081_/X hold704/X _2894_/S vssd1 vssd1 vccd1 vccd1 _2894_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1845_ _1845_/A _1871_/A _1871_/B vssd1 vssd1 vccd1 vccd1 _1846_/A sky130_fd_sc_hd__and3_1
XFILLER_0_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold602 _3470_/Q vssd1 vssd1 vccd1 vccd1 hold602/X sky130_fd_sc_hd__dlygate4sd3_1
X_1776_ _3626_/Q _3625_/Q vssd1 vssd1 vccd1 vccd1 _2056_/A sky130_fd_sc_hd__or2_4
Xhold624 _3339_/Q vssd1 vssd1 vccd1 vccd1 hold624/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold613 _2896_/X vssd1 vssd1 vccd1 vccd1 _3419_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 _2853_/X vssd1 vssd1 vccd1 vccd1 _3376_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3515_ _3614_/CLK _3515_/D _3009_/Y vssd1 vssd1 vccd1 vccd1 _3515_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold646 _3413_/Q vssd1 vssd1 vccd1 vccd1 hold646/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 _3181_/Q vssd1 vssd1 vccd1 vccd1 hold668/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 _2629_/X vssd1 vssd1 vccd1 vccd1 _3169_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 _2902_/X vssd1 vssd1 vccd1 vccd1 _3425_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3446_ _3636_/CLK _3446_/D _2940_/Y vssd1 vssd1 vccd1 vccd1 _3446_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ _3604_/CLK _3377_/D _2925_/Y vssd1 vssd1 vccd1 vccd1 _3377_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2328_ _3443_/Q _1601_/Y _2156_/B _2327_/X vssd1 vssd1 vccd1 vccd1 _2328_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_79_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2259_ _3467_/Q hold826/X _3466_/Q vssd1 vssd1 vccd1 vccd1 _2259_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_34_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3559_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2759__A1 _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1630_ _2393_/A hold7/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__nor2_1
X_1561_ _3635_/Q vssd1 vssd1 vccd1 vccd1 _2571_/A sky130_fd_sc_hd__inv_2
X_3300_ _3318_/CLK _3300_/D vssd1 vssd1 vccd1 vccd1 _3300_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _3612_/CLK _3231_/D vssd1 vssd1 vccd1 vccd1 _3231_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ _3404_/CLK _3162_/D vssd1 vssd1 vccd1 vccd1 _3162_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2695__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2113_ _2115_/A hold80/X vssd1 vssd1 vccd1 vccd1 _2114_/C sky130_fd_sc_hd__and2_1
X_3093_ _3124_/A vssd1 vssd1 vccd1 vccd1 _3093_/Y sky130_fd_sc_hd__inv_2
X_2044_ _3215_/Q _3206_/Q _3197_/Q _3323_/Q _2044_/S0 _2044_/S1 vssd1 vssd1 vccd1
+ vccd1 _2044_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_55_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2542__S0 _1943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2946_ _3128_/A vssd1 vssd1 vccd1 vccd1 _2946_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2877_ _2097_/A hold606/X _2884_/S vssd1 vssd1 vccd1 vccd1 _2877_/X sky130_fd_sc_hd__mux2_1
X_1828_ hold874/X hold861/X _1833_/S vssd1 vssd1 vccd1 vccd1 _3548_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_32_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold410 _3237_/Q vssd1 vssd1 vccd1 vccd1 hold410/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 _2733_/X vssd1 vssd1 vccd1 vccd1 _3259_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 _3212_/Q vssd1 vssd1 vccd1 vccd1 hold432/X sky130_fd_sc_hd__dlygate4sd3_1
X_1759_ _1811_/A _3564_/Q _1772_/B vssd1 vssd1 vccd1 vccd1 _1759_/X sky130_fd_sc_hd__or3_1
Xhold421 _2719_/X vssd1 vssd1 vccd1 vccd1 _3246_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 _3494_/Q vssd1 vssd1 vccd1 vccd1 hold454/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 _3483_/Q vssd1 vssd1 vccd1 vccd1 _2220_/S sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 _3482_/Q vssd1 vssd1 vccd1 vccd1 hold476/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 _3492_/Q vssd1 vssd1 vccd1 vccd1 _2179_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold498 _2198_/X vssd1 vssd1 vccd1 vccd1 _3488_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3429_ _3435_/CLK _3429_/D vssd1 vssd1 vccd1 vccd1 _3429_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2686__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2610__A0 _2342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1652__A1 hold86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2800_ hold402/X _2810_/A1 _2803_/S vssd1 vssd1 vccd1 vccd1 _2800_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2601__A0 _2097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2731_ _2811_/A1 hold416/X _2733_/S vssd1 vssd1 vccd1 vccd1 _2731_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_81_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2662_ _2794_/A _2794_/B vssd1 vssd1 vccd1 vccd1 _2804_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2593_ hold406/X _2809_/A1 _2597_/S vssd1 vssd1 vccd1 vccd1 _2593_/X sky130_fd_sc_hd__mux2_1
X_1613_ hold93/A _1613_/B _1625_/B hold17/X vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__or4_1
XFILLER_0_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2668__A0 _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3214_ _3513_/CLK _3214_/D vssd1 vssd1 vccd1 vccd1 _3214_/Q sky130_fd_sc_hd__dfxtp_1
X_3145_ _3414_/CLK _3145_/D vssd1 vssd1 vccd1 vccd1 _3145_/Q sky130_fd_sc_hd__dfxtp_1
X_3076_ _3124_/A vssd1 vssd1 vccd1 vccd1 _3076_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_82_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2515__S0 _1943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2027_ _1985_/S _2027_/B vssd1 vssd1 vccd1 vccd1 _2027_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2840__A0 _2079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1643__A1 _2395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2929_ _3128_/A vssd1 vssd1 vccd1 vccd1 _2929_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold251 _2777_/X vssd1 vssd1 vccd1 vccd1 _3298_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 _2664_/X vssd1 vssd1 vccd1 vccd1 _3197_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _2674_/X vssd1 vssd1 vccd1 vccd1 _3206_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 _2802_/X vssd1 vssd1 vccd1 vccd1 _3321_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 _3233_/Q vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _2727_/X vssd1 vssd1 vccd1 vccd1 _3253_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1643__S hold8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2659__A0 _2338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput8 input8/A vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_0__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_5_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2050__A1 _1985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2714_ _2794_/A _2794_/B _2764_/A vssd1 vssd1 vccd1 vccd1 _2723_/S sky130_fd_sc_hd__or3_4
X_2645_ _2105_/B hold692/X _2650_/S vssd1 vssd1 vccd1 vccd1 _2645_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2889__A0 _2104_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2576_ _2583_/B _2576_/B vssd1 vssd1 vccd1 vccd1 _2576_/X sky130_fd_sc_hd__and2_2
X_3128_ _3128_/A vssd1 vssd1 vccd1 vccd1 _3128_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_69_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3059_ _3065_/A vssd1 vssd1 vccd1 vccd1 _3059_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1638__S hold8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2041__A1 _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2993__A _3131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2430_ _2429_/X _2428_/X _2551_/S vssd1 vssd1 vccd1 vccd1 _2430_/X sky130_fd_sc_hd__mux2_1
X_2361_ _3563_/Q _3562_/Q _3561_/Q _3560_/Q vssd1 vssd1 vccd1 vccd1 _2361_/X sky130_fd_sc_hd__or4_1
XANTENNA__3064__A _3131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2292_ _3459_/Q hold83/X hold30/X vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__mux2_1
XFILLER_0_2_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout124_A _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2628_ _2338_/B hold796/X _2629_/S vssd1 vssd1 vccd1 vccd1 _2628_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2559_ _3623_/Q _1645_/Y _2493_/Y _2557_/X _2558_/X vssd1 vssd1 vccd1 vccd1 _2559_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2752__S _2753_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2262__A1 _2231_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1999__S1 _2044_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1930_ _1930_/A _1930_/B vssd1 vssd1 vccd1 vccd1 _1930_/X sky130_fd_sc_hd__and2_1
XFILLER_0_56_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1861_ _1583_/A _1850_/A _1835_/A vssd1 vssd1 vccd1 vccd1 _1861_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_56_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3600_ _3604_/CLK _3600_/D _3091_/Y vssd1 vssd1 vccd1 vccd1 _3600_/Q sky130_fd_sc_hd__dfrtp_1
Xinput22 hold40/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__clkbuf_2
Xinput11 hold4/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__buf_1
X_3531_ _3539_/CLK _3531_/D _3025_/Y vssd1 vssd1 vccd1 vccd1 _3531_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1792_ _2383_/C _1792_/B _1792_/C vssd1 vssd1 vccd1 vccd1 _1793_/A sky130_fd_sc_hd__and3_1
Xinput33 hold43/X vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold817 _1998_/X vssd1 vssd1 vccd1 vccd1 _3510_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 _3505_/Q vssd1 vssd1 vccd1 vccd1 hold828/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold806 _3589_/Q vssd1 vssd1 vccd1 vccd1 hold806/X sky130_fd_sc_hd__dlygate4sd3_1
X_3462_ _3637_/CLK _3462_/D _2956_/Y vssd1 vssd1 vccd1 vccd1 _3462_/Q sky130_fd_sc_hd__dfrtp_1
Xhold839 _1697_/X vssd1 vssd1 vccd1 vccd1 _3579_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2413_ _3596_/Q _2568_/B _2441_/B vssd1 vssd1 vccd1 vccd1 _2413_/X sky130_fd_sc_hd__o21ba_1
X_3393_ _3423_/CLK _3393_/D vssd1 vssd1 vccd1 vccd1 _3393_/Q sky130_fd_sc_hd__dfxtp_1
X_2344_ _2344_/A _2344_/B _2344_/C _2344_/D vssd1 vssd1 vccd1 vccd1 _2344_/X sky130_fd_sc_hd__and4_1
X_2275_ _2275_/A _2278_/B vssd1 vssd1 vccd1 vccd1 _2275_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__2492__A1 _3341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2747__S _2753_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xuart_macro_wrapper_135 vssd1 vssd1 vccd1 vccd1 uart_macro_wrapper_135/HI wbs_dat_o[24]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3523_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2016__A_N _1985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2060_ _3549_/Q _2089_/B vssd1 vssd1 vccd1 vccd1 _2060_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2962_ _3044_/A vssd1 vssd1 vccd1 vccd1 _2962_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1913_ _1912_/A _1910_/B _1910_/Y _2163_/B vssd1 vssd1 vccd1 vccd1 _3522_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2893_ _2076_/X hold740/X _2894_/S vssd1 vssd1 vccd1 vccd1 _2893_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1844_ _1871_/A _1871_/B vssd1 vssd1 vccd1 vccd1 _1844_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold603 _2251_/X vssd1 vssd1 vccd1 vccd1 _3475_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1775_ _1795_/B _1775_/B vssd1 vssd1 vccd1 vccd1 _1775_/Y sky130_fd_sc_hd__nand2_1
Xhold614 _3191_/Q vssd1 vssd1 vccd1 vccd1 hold614/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 _2822_/X vssd1 vssd1 vccd1 vccd1 _3339_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold636 _3412_/Q vssd1 vssd1 vccd1 vccd1 hold636/X sky130_fd_sc_hd__dlygate4sd3_1
X_3514_ _3623_/CLK _3514_/D _3008_/Y vssd1 vssd1 vccd1 vccd1 _3514_/Q sky130_fd_sc_hd__dfrtp_1
X_3445_ _3540_/CLK _3445_/D _2939_/Y vssd1 vssd1 vccd1 vccd1 _3445_/Q sky130_fd_sc_hd__dfrtp_1
Xhold647 _2889_/X vssd1 vssd1 vccd1 vccd1 _3413_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold669 _2644_/X vssd1 vssd1 vccd1 vccd1 _3181_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 _3416_/Q vssd1 vssd1 vccd1 vccd1 hold658/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _3427_/CLK _3376_/D vssd1 vssd1 vccd1 vccd1 _3376_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2327_ hold828/X _3346_/Q _1956_/B _2145_/A _3345_/Q vssd1 vssd1 vccd1 vccd1 _2327_/X
+ sky130_fd_sc_hd__a2111o_1
X_2258_ hold917/X hold922/X _2258_/S vssd1 vssd1 vccd1 vccd1 _3468_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2189_ _2214_/A _2196_/B vssd1 vssd1 vccd1 vccd1 _2189_/X sky130_fd_sc_hd__or2_1
XFILLER_0_62_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2000__S0 _2044_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1560_ _1834_/A vssd1 vssd1 vccd1 vccd1 _1560_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_1_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _3612_/CLK _3230_/D vssd1 vssd1 vccd1 vccd1 _3230_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ _3526_/CLK _3161_/D vssd1 vssd1 vccd1 vccd1 _3161_/Q sky130_fd_sc_hd__dfxtp_1
X_2112_ _2112_/A _2112_/B vssd1 vssd1 vccd1 vccd1 _2116_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3092_ _3095_/A vssd1 vssd1 vccd1 vccd1 _3092_/Y sky130_fd_sc_hd__inv_2
X_2043_ hold307/X hold360/X hold284/X hold282/X _2044_/S0 _2044_/S1 vssd1 vssd1 vccd1
+ vccd1 _2043_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2542__S1 _2550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2945_ _3128_/A vssd1 vssd1 vccd1 vccd1 _2945_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2876_ _2342_/B hold582/X _2884_/S vssd1 vssd1 vccd1 vccd1 _2876_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1827_ hold830/X _3549_/Q _1831_/S vssd1 vssd1 vccd1 vccd1 _1827_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold411 _2709_/X vssd1 vssd1 vccd1 vccd1 _3237_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold400 _3228_/Q vssd1 vssd1 vccd1 vccd1 hold400/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 _3446_/Q vssd1 vssd1 vccd1 vccd1 hold444/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold433 _2680_/X vssd1 vssd1 vccd1 vccd1 _3212_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1758_ hold973/X _2383_/C _1757_/X vssd1 vssd1 vccd1 vccd1 _1758_/X sky130_fd_sc_hd__o21a_1
Xhold422 _3264_/Q vssd1 vssd1 vccd1 vccd1 hold422/X sky130_fd_sc_hd__dlygate4sd3_1
X_1689_ hold241/X _2395_/A hold21/X vssd1 vssd1 vccd1 vccd1 _3597_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_40_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold466 _2178_/X vssd1 vssd1 vccd1 vccd1 _2180_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 _2245_/X vssd1 vssd1 vccd1 vccd1 hold455/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 _2230_/X vssd1 vssd1 vccd1 vccd1 _3482_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 _2220_/X vssd1 vssd1 vccd1 vccd1 _3483_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3428_ _3523_/CLK _3428_/D vssd1 vssd1 vccd1 vccd1 _3428_/Q sky130_fd_sc_hd__dfxtp_1
Xhold499 hold499/A vssd1 vssd1 vccd1 vccd1 _1940_/S sky130_fd_sc_hd__buf_1
XANTENNA__2297__S hold30/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3359_ _3403_/CLK _3359_/D vssd1 vssd1 vccd1 vccd1 _3359_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2760__S _2763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2677__A1 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2670__S _2672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2730_ _2810_/A1 hold335/X _2733_/S vssd1 vssd1 vccd1 vccd1 _2730_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2661_ _3491_/Q _2661_/B _3492_/Q vssd1 vssd1 vccd1 vccd1 _2784_/C sky130_fd_sc_hd__nand3b_2
X_1612_ hold27/X _1612_/B vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__nor2_2
X_2592_ hold136/X _2808_/A1 _2594_/S vssd1 vssd1 vccd1 vccd1 _2592_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3213_ _3330_/CLK _3213_/D vssd1 vssd1 vccd1 vccd1 _3213_/Q sky130_fd_sc_hd__dfxtp_1
X_3144_ _3435_/CLK _3144_/D vssd1 vssd1 vccd1 vccd1 _3144_/Q sky130_fd_sc_hd__dfxtp_1
X_3075_ _3126_/A vssd1 vssd1 vccd1 vccd1 _3075_/Y sky130_fd_sc_hd__inv_2
X_2026_ _2025_/X _2024_/X _2045_/S vssd1 vssd1 vccd1 vccd1 _2027_/B sky130_fd_sc_hd__mux2_1
XANTENNA__2515__S1 _2550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2928_ _3095_/A vssd1 vssd1 vccd1 vccd1 _2928_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_72_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2859_ _2105_/B hold726/X _2864_/S vssd1 vssd1 vccd1 vccd1 _2859_/X sky130_fd_sc_hd__mux2_1
Xhold252 _3260_/Q vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 _3597_/Q vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2451__S0 _2554_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold230 _2687_/X vssd1 vssd1 vccd1 vccd1 _3217_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 _3269_/Q vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 _3249_/Q vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 _2705_/X vssd1 vssd1 vccd1 vccd1 _3233_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _3136_/Q vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2755__S _2763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2831__A1 _2075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2490__S _3522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2665__S _2672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_59_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2822__A1 _2338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2713_ _2813_/A1 hold436/X _2713_/S vssd1 vssd1 vccd1 vccd1 _2713_/X sky130_fd_sc_hd__mux2_1
X_2644_ _2105_/A hold668/X _2650_/S vssd1 vssd1 vccd1 vccd1 _2644_/X sky130_fd_sc_hd__mux2_1
X_2575_ _2511_/Y _2581_/C _2574_/X _2511_/B _3456_/Q vssd1 vssd1 vccd1 vccd1 _2576_/B
+ sky130_fd_sc_hd__a32o_1
X_3127_ _3128_/A vssd1 vssd1 vccd1 vccd1 _3127_/Y sky130_fd_sc_hd__inv_2
X_3058_ _3121_/A vssd1 vssd1 vccd1 vccd1 _3058_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2813__A1 _2813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2009_ hold824/X _2008_/X _2053_/S vssd1 vssd1 vccd1 vccd1 _2009_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2041__A2 _2039_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold114_A _2287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2740__A0 _2810_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2360_ _1597_/Y _2359_/X hold512/X vssd1 vssd1 vccd1 vccd1 _2360_/Y sky130_fd_sc_hd__a21oi_1
X_2291_ _2393_/A hold29/X vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__nor2_2
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2627_ _2075_/B hold666/X _2629_/S vssd1 vssd1 vccd1 vccd1 _2627_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_28_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3580_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2731__A0 _2811_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2558_ _3380_/Q _1678_/X _2412_/Y hold74/A vssd1 vssd1 vccd1 vccd1 _2558_/X sky130_fd_sc_hd__o211a_1
X_2489_ _2488_/X _2487_/X _3521_/Q vssd1 vssd1 vccd1 vccd1 _2489_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_65_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2722__A0 _2812_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2789__A0 _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1860_ _1835_/A _1852_/Y _1859_/X _1859_/A _1560_/Y vssd1 vssd1 vccd1 vccd1 _1860_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_56_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput12 input12/A vssd1 vssd1 vccd1 vccd1 _1624_/C sky130_fd_sc_hd__clkbuf_2
X_1791_ _1791_/A _1791_/B _2123_/A _1791_/D vssd1 vssd1 vccd1 vccd1 _1792_/C sky130_fd_sc_hd__and4_1
X_3530_ _3539_/CLK _3530_/D _3024_/Y vssd1 vssd1 vccd1 vccd1 _3530_/Q sky130_fd_sc_hd__dfrtp_1
Xinput34 hold48/X vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__buf_1
Xinput23 hold75/X vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold818 hold818/A vssd1 vssd1 vccd1 vccd1 _1711_/B sky130_fd_sc_hd__buf_1
Xhold807 _2349_/X vssd1 vssd1 vccd1 vccd1 _3377_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3461_ _3637_/CLK _3461_/D _2955_/Y vssd1 vssd1 vccd1 vccd1 _3461_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3075__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold829 _2053_/X vssd1 vssd1 vccd1 vccd1 _3505_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3392_ _3523_/CLK _3392_/D vssd1 vssd1 vccd1 vccd1 _3392_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2713__A0 _2813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2412_ hold20/A _2416_/A vssd1 vssd1 vccd1 vccd1 _2412_/Y sky130_fd_sc_hd__nand2_1
X_2343_ _1571_/Y _2105_/A _2338_/Y _2339_/Y _1889_/Y vssd1 vssd1 vccd1 vccd1 _2344_/D
+ sky130_fd_sc_hd__o2111a_1
X_2274_ _2277_/A _2280_/B vssd1 vssd1 vccd1 vccd1 _2278_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1989_ hold302/X hold321/X hold323/X hold351/X _2044_/S0 _2044_/S1 vssd1 vssd1 vccd1
+ vccd1 _1989_/X sky130_fd_sc_hd__mux4_1
X_3659_ _3659_/A vssd1 vssd1 vccd1 vccd1 _3659_/X sky130_fd_sc_hd__buf_1
XFILLER_0_2_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2763__S _2763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire80 wire80/A vssd1 vssd1 vccd1 vccd1 wire80/X sky130_fd_sc_hd__buf_1
XFILLER_0_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xuart_macro_wrapper_136 vssd1 vssd1 vccd1 vccd1 uart_macro_wrapper_136/HI wbs_dat_o[29]
+ sky130_fd_sc_hd__conb_1
XFILLER_0_80_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_2_3__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2961_ _3044_/A vssd1 vssd1 vccd1 vccd1 _2961_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_56_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1912_ _1912_/A _1915_/A vssd1 vssd1 vccd1 vccd1 _2163_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_29_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2892_ _2074_/X hold658/X _2894_/S vssd1 vssd1 vccd1 vccd1 _2892_/X sky130_fd_sc_hd__mux2_1
X_1843_ _1843_/A _1843_/B vssd1 vssd1 vccd1 vccd1 _1871_/B sky130_fd_sc_hd__and2_1
XFILLER_0_44_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1774_ _1745_/B _1744_/A _1774_/C _3552_/Q vssd1 vssd1 vccd1 vccd1 _1775_/B sky130_fd_sc_hd__and4bb_1
Xhold615 _2655_/X vssd1 vssd1 vccd1 vccd1 _3191_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 _3431_/Q vssd1 vssd1 vccd1 vccd1 hold626/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold604 _3434_/Q vssd1 vssd1 vccd1 vccd1 hold604/X sky130_fd_sc_hd__dlygate4sd3_1
X_3513_ _3513_/CLK _3513_/D _3007_/Y vssd1 vssd1 vccd1 vccd1 _3513_/Q sky130_fd_sc_hd__dfrtp_1
X_3444_ _3540_/CLK _3444_/D _2938_/Y vssd1 vssd1 vccd1 vccd1 _3444_/Q sky130_fd_sc_hd__dfrtp_1
Xhold637 _2888_/X vssd1 vssd1 vccd1 vccd1 _3412_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold659 _2892_/X vssd1 vssd1 vccd1 vccd1 _3416_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 _3158_/Q vssd1 vssd1 vccd1 vccd1 hold648/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ _3583_/CLK _3375_/D vssd1 vssd1 vccd1 vccd1 _3375_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2326_ _2114_/C _2115_/Y _2326_/S vssd1 vssd1 vccd1 vccd1 _2326_/X sky130_fd_sc_hd__mux2_1
X_2257_ hold853/X hold917/X _2258_/S vssd1 vssd1 vccd1 vccd1 _3469_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1673__A0 _2396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2188_ _2214_/A _2185_/Y _2202_/A vssd1 vssd1 vccd1 vccd1 _2188_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_43_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3526_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout97_A _2224_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2758__S _2763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2000__S1 _2044_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2668__S _2672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _3427_/CLK _3160_/D vssd1 vssd1 vccd1 vccd1 _3160_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
X_3091_ _3095_/A vssd1 vssd1 vccd1 vccd1 _3091_/Y sky130_fd_sc_hd__inv_2
X_2111_ _2111_/A _2111_/B vssd1 vssd1 vccd1 vccd1 _2112_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2042_ hold820/X _2041_/Y _2053_/S vssd1 vssd1 vccd1 vccd1 _2042_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2944_ _3133_/A vssd1 vssd1 vccd1 vccd1 _2944_/Y sky130_fd_sc_hd__inv_2
X_2875_ _2875_/A _2875_/B vssd1 vssd1 vccd1 vccd1 _2884_/S sky130_fd_sc_hd__or2_4
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1826_ hold855/X hold830/X _1831_/S vssd1 vssd1 vccd1 vccd1 _1826_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2907__A0 _2097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold401 _2699_/X vssd1 vssd1 vccd1 vccd1 _3228_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 _3293_/Q vssd1 vssd1 vccd1 vccd1 hold434/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 _3329_/Q vssd1 vssd1 vccd1 vccd1 hold412/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 _3140_/Q vssd1 vssd1 vccd1 vccd1 hold445/X sky130_fd_sc_hd__dlygate4sd3_1
X_1757_ _1811_/A _3565_/Q _1772_/B vssd1 vssd1 vccd1 vccd1 _1757_/X sky130_fd_sc_hd__or3_1
Xhold423 _2739_/X vssd1 vssd1 vccd1 vccd1 _3264_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1688_ hold304/X _2396_/A hold21/X vssd1 vssd1 vccd1 vccd1 _3598_/D sky130_fd_sc_hd__mux2_1
Xhold478 hold478/A vssd1 vssd1 vccd1 vccd1 _3583_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 _2180_/X vssd1 vssd1 vccd1 vccd1 _3492_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 _2246_/X vssd1 vssd1 vccd1 vccd1 _3476_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3427_ _3427_/CLK _3427_/D vssd1 vssd1 vccd1 vccd1 _3427_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2135__A1 _2052_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold489 _3516_/Q vssd1 vssd1 vccd1 vccd1 _2350_/B sky130_fd_sc_hd__clkbuf_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ _3427_/CLK _3358_/D vssd1 vssd1 vccd1 vccd1 _3358_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _1565_/Y _2056_/B _1996_/A vssd1 vssd1 vccd1 vccd1 _2310_/B sky130_fd_sc_hd__a21oi_1
X_3289_ _3316_/CLK _3289_/D vssd1 vssd1 vccd1 vccd1 _3289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold990 _2154_/X vssd1 vssd1 vccd1 vccd1 _3499_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1980__S0 _2224_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2660_ _2339_/B hold730/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2660_/X sky130_fd_sc_hd__mux2_1
X_1611_ _1660_/A hold65/A input4/X input5/X vssd1 vssd1 vccd1 vccd1 _1611_/X sky130_fd_sc_hd__or4_1
X_2591_ hold274/X _2807_/A1 _2594_/S vssd1 vssd1 vccd1 vccd1 _2591_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3212_ _3331_/CLK _3212_/D vssd1 vssd1 vccd1 vccd1 _3212_/Q sky130_fd_sc_hd__dfxtp_1
X_3143_ _3403_/CLK _3143_/D vssd1 vssd1 vccd1 vccd1 _3143_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1971__S0 _1590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3074_ _3114_/A vssd1 vssd1 vccd1 vccd1 _3074_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_82_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2025_ _3244_/Q _3316_/Q _3307_/Q _3298_/Q _1590_/A _2222_/A vssd1 vssd1 vccd1 vccd1
+ _2025_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2861__S _2864_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2927_ _3133_/A vssd1 vssd1 vccd1 vccd1 _2927_/Y sky130_fd_sc_hd__inv_2
X_2858_ _2105_/A hold800/X _2864_/S vssd1 vssd1 vccd1 vccd1 _2858_/X sky130_fd_sc_hd__mux2_1
Xhold220 _2767_/X vssd1 vssd1 vccd1 vccd1 _3289_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1809_ _1815_/B _1809_/B vssd1 vssd1 vccd1 vccd1 _1810_/A sky130_fd_sc_hd__nor2_1
X_2789_ _2809_/A1 hold438/X _2793_/S vssd1 vssd1 vccd1 vccd1 _2789_/X sky130_fd_sc_hd__mux2_1
Xhold231 _3262_/Q vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 _2735_/X vssd1 vssd1 vccd1 vccd1 _3260_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2451__S1 _1911_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold242 _3215_/Q vssd1 vssd1 vccd1 vccd1 hold242/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _2745_/X vssd1 vssd1 vccd1 vccd1 _3269_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold286 _3323_/Q vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 _2591_/X vssd1 vssd1 vccd1 vccd1 _3136_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 _2722_/X vssd1 vssd1 vccd1 vccd1 _3249_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1962__S0 _1590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1619__A0 _3642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2771__S _2773_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2595__A1 _2811_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2681__S _2682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2712_ _2812_/A1 hold396/X _2713_/S vssd1 vssd1 vccd1 vccd1 _2712_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2643_ _2097_/A hold654/X _2650_/S vssd1 vssd1 vccd1 vccd1 _2643_/X sky130_fd_sc_hd__mux2_1
X_2574_ _3636_/Q hold7/A vssd1 vssd1 vccd1 vccd1 _2574_/X sky130_fd_sc_hd__or2_1
XFILLER_0_10_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2856__S _2864_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3126_ _3126_/A vssd1 vssd1 vccd1 vccd1 _3126_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3057_ _3121_/A vssd1 vssd1 vccd1 vccd1 _3057_/Y sky130_fd_sc_hd__inv_2
X_2008_ hold816/X _2007_/Y _2052_/S vssd1 vssd1 vccd1 vccd1 _2008_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1996__A _1996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2766__S _2773_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output60_A _3659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2290_ hold28/X _2419_/B vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__nand2_4
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2676__S _2682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2626_ _2079_/A hold780/X _2629_/S vssd1 vssd1 vccd1 vccd1 _2626_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2557_ _3380_/Q _3592_/Q _2568_/C vssd1 vssd1 vccd1 vccd1 _2557_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2488_ _3173_/Q _3422_/Q _3413_/Q _3155_/Q _2554_/S0 _1911_/B vssd1 vssd1 vccd1 vccd1
+ _2488_/X sky130_fd_sc_hd__mux4_1
X_3109_ _3114_/A vssd1 vssd1 vccd1 vccd1 _3109_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2798__A1 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 input13/A vssd1 vssd1 vccd1 vccd1 _1613_/B sky130_fd_sc_hd__buf_1
XFILLER_0_24_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1790_ _3557_/Q _2124_/B _1786_/Y _1787_/X vssd1 vssd1 vccd1 vccd1 _1791_/D sky130_fd_sc_hd__o211a_1
Xinput24 hold35/X vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__buf_1
Xinput35 hold13/X vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold819 _1711_/X vssd1 vssd1 vccd1 vccd1 _3572_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold808 _3511_/Q vssd1 vssd1 vccd1 vccd1 hold808/X sky130_fd_sc_hd__dlygate4sd3_1
X_3460_ _3637_/CLK _3460_/D _2954_/Y vssd1 vssd1 vccd1 vccd1 _3460_/Q sky130_fd_sc_hd__dfrtp_1
X_3391_ _3436_/CLK _3391_/D vssd1 vssd1 vccd1 vccd1 _3391_/Q sky130_fd_sc_hd__dfxtp_1
X_2411_ hold20/A _2416_/A vssd1 vssd1 vccd1 vccd1 _2568_/B sky130_fd_sc_hd__and2_2
XFILLER_0_20_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2342_ _2342_/A _2342_/B vssd1 vssd1 vccd1 vccd1 _2344_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2273_ _2273_/A _2273_/B _2283_/B vssd1 vssd1 vccd1 vccd1 _2280_/B sky130_fd_sc_hd__and3_1
XFILLER_0_47_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1988_ hold335/X hold430/X hold315/X hold311/X _2044_/S0 _2044_/S1 vssd1 vssd1 vccd1
+ vccd1 _1988_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3658_ _3659_/A vssd1 vssd1 vccd1 vccd1 _3658_/X sky130_fd_sc_hd__buf_1
X_2609_ _3526_/Q _2905_/B _2905_/C vssd1 vssd1 vccd1 vccd1 _2618_/S sky130_fd_sc_hd__or3b_4
X_3589_ _3614_/CLK hold34/X _3080_/Y vssd1 vssd1 vccd1 vccd1 _3589_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2640__A0 _2339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xuart_macro_wrapper_137 vssd1 vssd1 vccd1 vccd1 io_oeb[0] uart_macro_wrapper_137/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_46_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_88_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2554__S0 _2554_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1682__A1 hold49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2960_ _3073_/A vssd1 vssd1 vccd1 vccd1 _2960_/Y sky130_fd_sc_hd__inv_2
X_2891_ _2067_/Y hold586/X _2894_/S vssd1 vssd1 vccd1 vccd1 _2891_/X sky130_fd_sc_hd__mux2_1
X_1911_ _1911_/A _1911_/B _1911_/C vssd1 vssd1 vccd1 vccd1 _1915_/A sky130_fd_sc_hd__and3_1
XFILLER_0_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1842_ _1843_/B vssd1 vssd1 vccd1 vccd1 _1842_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1773_ _1767_/B _2383_/C _1772_/X vssd1 vssd1 vccd1 vccd1 _1773_/X sky130_fd_sc_hd__o21a_1
Xhold627 _2909_/X vssd1 vssd1 vccd1 vccd1 _3431_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 _3426_/Q vssd1 vssd1 vccd1 vccd1 hold616/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold605 _2912_/X vssd1 vssd1 vccd1 vccd1 _3434_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3512_ _3612_/CLK _3512_/D _3006_/Y vssd1 vssd1 vccd1 vccd1 _3512_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold638 _3364_/Q vssd1 vssd1 vccd1 vccd1 hold638/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 _2616_/X vssd1 vssd1 vccd1 vccd1 _3158_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3443_ _3580_/CLK _3443_/D _2937_/Y vssd1 vssd1 vccd1 vccd1 _3443_/Q sky130_fd_sc_hd__dfstp_2
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2698__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _3416_/CLK _3374_/D vssd1 vssd1 vccd1 vccd1 _3374_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2325_ _2314_/Y _2323_/Y _2324_/Y vssd1 vssd1 vccd1 vccd1 _2326_/S sky130_fd_sc_hd__o21a_1
X_2256_ hold602/X hold853/X _3466_/Q vssd1 vssd1 vccd1 vccd1 _2256_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2545__S0 _2554_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2864__S _2864_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2187_ _2187_/A _2214_/A _2661_/B _2200_/B vssd1 vssd1 vccd1 vccd1 _2202_/A sky130_fd_sc_hd__or4_1
XANTENNA__2622__A0 _2097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_12_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3305_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2689__A0 _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2861__A0 _2079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1664__A1 _2397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2613__A0 _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
X_2110_ _2111_/B vssd1 vssd1 vccd1 vccd1 _2110_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_55_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3090_ _3095_/A vssd1 vssd1 vccd1 vccd1 _3090_/Y sky130_fd_sc_hd__inv_2
X_2041_ _3346_/Q _2039_/Y _2040_/Y vssd1 vssd1 vccd1 vccd1 _2041_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2852__A0 _2338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1655__A1 _2395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2943_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2943_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2604__A0 _2111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2874_ hold518/X _2339_/B _2874_/S vssd1 vssd1 vccd1 vccd1 _2874_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1825_ _2111_/A hold855/X _1833_/S vssd1 vssd1 vccd1 vccd1 _1825_/X sky130_fd_sc_hd__mux2_1
Xhold402 _3319_/Q vssd1 vssd1 vccd1 vccd1 hold402/X sky130_fd_sc_hd__dlygate4sd3_1
X_1756_ hold967/X _2383_/C _1755_/X vssd1 vssd1 vccd1 vccd1 _1756_/X sky130_fd_sc_hd__o21a_1
Xhold435 _2771_/X vssd1 vssd1 vccd1 vccd1 _3293_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2859__S _2864_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold413 _2811_/X vssd1 vssd1 vccd1 vccd1 _3329_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 _3318_/Q vssd1 vssd1 vccd1 vccd1 hold424/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 _3223_/Q vssd1 vssd1 vccd1 vccd1 hold457/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 hold468/A vssd1 vssd1 vccd1 vccd1 _1933_/A sky130_fd_sc_hd__clkbuf_4
Xhold446 _2595_/X vssd1 vssd1 vccd1 vccd1 _3140_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1687_ hold201/X _2397_/A hold21/X vssd1 vssd1 vccd1 vccd1 _3599_/D sky130_fd_sc_hd__mux2_1
X_3426_ _3583_/CLK _3426_/D vssd1 vssd1 vccd1 vccd1 _3426_/Q sky130_fd_sc_hd__dfxtp_1
Xhold479 _3514_/Q vssd1 vssd1 vccd1 vccd1 _1891_/A sky130_fd_sc_hd__buf_2
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3357_ _3369_/CLK _3357_/D vssd1 vssd1 vccd1 vccd1 _3357_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _1565_/Y _1780_/Y _2007_/A vssd1 vssd1 vccd1 vccd1 _2310_/A sky130_fd_sc_hd__a21oi_1
X_3288_ _3319_/CLK _3288_/D vssd1 vssd1 vccd1 vccd1 _3288_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2518__S0 _2554_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2239_ _2260_/B _2241_/A vssd1 vssd1 vccd1 vccd1 _2239_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_67_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2843__A0 _2339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2342__B _2342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2769__S _2773_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold991 _3536_/Q vssd1 vssd1 vccd1 vccd1 _1584_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold980 _1806_/Y vssd1 vssd1 vccd1 vccd1 _1807_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1980__S1 _2193_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1637__A1 hold44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2009__S _2053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1610_ input6/X input7/X hold26/X input9/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__or4_1
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2590_ hold202/X _2806_/A1 _2594_/S vssd1 vssd1 vccd1 vccd1 _2590_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2679__S _2682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3211_ _3328_/CLK _3211_/D vssd1 vssd1 vccd1 vccd1 _3211_/Q sky130_fd_sc_hd__dfxtp_1
X_3142_ _3513_/CLK _3142_/D vssd1 vssd1 vccd1 vccd1 _3142_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1971__S1 _2193_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3073_ _3073_/A vssd1 vssd1 vccd1 vccd1 _3073_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_82_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2024_ _3289_/Q _3280_/Q _3271_/Q _3262_/Q _1590_/A _2222_/A vssd1 vssd1 vccd1 vccd1
+ _2024_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_49_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2926_ _3133_/A vssd1 vssd1 vccd1 vccd1 _2926_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2857_ _2097_/A hold756/X _2864_/S vssd1 vssd1 vccd1 vccd1 _2857_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1808_ _1808_/A _1808_/B _1824_/A _1808_/D vssd1 vssd1 vccd1 vccd1 _1809_/B sky130_fd_sc_hd__or4_1
Xhold210 _3595_/Q vssd1 vssd1 vccd1 vccd1 _2214_/A sky130_fd_sc_hd__clkbuf_4
X_2788_ _2808_/A1 hold163/X _2793_/S vssd1 vssd1 vccd1 vccd1 _2788_/X sky130_fd_sc_hd__mux2_1
Xhold232 _2737_/X vssd1 vssd1 vccd1 vccd1 _3262_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 _3296_/Q vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
X_1739_ _1851_/A _3456_/Q _1726_/X _1728_/X _1731_/X vssd1 vssd1 vccd1 vccd1 _1741_/C
+ sky130_fd_sc_hd__a2111o_1
Xhold243 _2685_/X vssd1 vssd1 vccd1 vccd1 _3215_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 _3312_/Q vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 _3287_/Q vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 _3596_/Q vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 _2805_/X vssd1 vssd1 vccd1 vccd1 _3323_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3409_ _3436_/CLK _3409_/D vssd1 vssd1 vccd1 vccd1 _3409_/Q sky130_fd_sc_hd__dfxtp_1
Xhold298 _3615_/Q vssd1 vssd1 vccd1 vccd1 _2342_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1962__S1 _2193_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1619__A1 hold86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2711_ _2811_/A1 hold426/X _2713_/S vssd1 vssd1 vccd1 vccd1 _2711_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2642_ _2342_/B hold690/X _2650_/S vssd1 vssd1 vccd1 vccd1 _2642_/X sky130_fd_sc_hd__mux2_1
X_2573_ _2583_/B _2573_/B vssd1 vssd1 vccd1 vccd1 _2573_/X sky130_fd_sc_hd__and2_2
XANTENNA__1607__A _1609_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold30_A hold30/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3125_ _3126_/A vssd1 vssd1 vccd1 vccd1 _3125_/Y sky130_fd_sc_hd__inv_2
X_3056_ _3121_/A vssd1 vssd1 vccd1 vccd1 _3056_/Y sky130_fd_sc_hd__inv_2
X_2007_ _2007_/A vssd1 vssd1 vccd1 vccd1 _2007_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_45_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2909_ _2105_/B hold626/X _2914_/S vssd1 vssd1 vccd1 vccd1 _2909_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2017__A1 _1985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2692__S _2693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3089__A _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2625_ _2111_/B hold720/X _2629_/S vssd1 vssd1 vccd1 vccd1 _2625_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2556_ _3522_/Q _2556_/B vssd1 vssd1 vccd1 vccd1 _2556_/X sky130_fd_sc_hd__or2_1
X_2487_ _3371_/Q _3353_/Q _3362_/Q _3191_/Q _2554_/S0 _1911_/B vssd1 vssd1 vccd1 vccd1
+ _2487_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3108_ _3114_/A vssd1 vssd1 vccd1 vccd1 _3108_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_37_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3583_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3039_ _3044_/A vssd1 vssd1 vccd1 vccd1 _3039_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput25 hold10/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__clkbuf_1
Xinput36 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _1609_/A sky130_fd_sc_hd__buf_2
Xinput14 hold92/X vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold809 _1987_/X vssd1 vssd1 vccd1 vccd1 _3511_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2410_ _2410_/A _2415_/A vssd1 vssd1 vccd1 vccd1 _2416_/A sky130_fd_sc_hd__nand2_1
X_3390_ _3435_/CLK _3390_/D vssd1 vssd1 vccd1 vccd1 _3390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2341_ _1569_/Y _2079_/A _2075_/B _1568_/Y vssd1 vssd1 vccd1 vccd1 _2344_/B sky130_fd_sc_hd__a22oi_1
XANTENNA__2687__S _2693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2272_ _2272_/A _2272_/B _2272_/C vssd1 vssd1 vccd1 vccd1 _2283_/B sky130_fd_sc_hd__and3_1
XANTENNA__2021__S0 _2044_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1987_ hold808/X _1986_/X _2053_/S vssd1 vssd1 vccd1 vccd1 _1987_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout122_A _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3657_ _3659_/A vssd1 vssd1 vccd1 vccd1 _3657_/X sky130_fd_sc_hd__buf_1
XFILLER_0_2_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2608_ _2339_/B hold628/X _2608_/S vssd1 vssd1 vccd1 vccd1 _2608_/X sky130_fd_sc_hd__mux2_1
X_3588_ _3604_/CLK _3588_/D _3079_/Y vssd1 vssd1 vccd1 vccd1 _3588_/Q sky130_fd_sc_hd__dfrtp_1
X_2539_ hold69/A _1645_/Y _2568_/D _2537_/X vssd1 vssd1 vccd1 vccd1 _2539_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_38_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2003__S0 _2224_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2554__S1 _1942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_84_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2890_ _2109_/X hold728/X _2894_/S vssd1 vssd1 vccd1 vccd1 _2890_/X sky130_fd_sc_hd__mux2_1
X_1910_ _1933_/A _1910_/B vssd1 vssd1 vccd1 vccd1 _1910_/Y sky130_fd_sc_hd__nor2_1
X_1841_ _1841_/A _1877_/A _1877_/B vssd1 vssd1 vccd1 vccd1 _1843_/B sky130_fd_sc_hd__and3_1
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1772_ _1811_/A _1772_/B _2111_/A vssd1 vssd1 vccd1 vccd1 _1772_/X sky130_fd_sc_hd__or3_1
Xhold606 _3402_/Q vssd1 vssd1 vccd1 vccd1 hold606/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 _2903_/X vssd1 vssd1 vccd1 vccd1 _3426_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3511_ _3612_/CLK _3511_/D _3005_/Y vssd1 vssd1 vccd1 vccd1 _3511_/Q sky130_fd_sc_hd__dfrtp_1
Xhold639 _2840_/X vssd1 vssd1 vccd1 vccd1 _3364_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 _3151_/Q vssd1 vssd1 vccd1 vccd1 hold628/X sky130_fd_sc_hd__dlygate4sd3_1
X_3442_ _3551_/CLK _3442_/D _2936_/Y vssd1 vssd1 vccd1 vccd1 _3442_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ _3416_/CLK _3373_/D vssd1 vssd1 vccd1 vccd1 _3373_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _2314_/Y _2323_/Y hold70/X vssd1 vssd1 vccd1 vccd1 _2324_/Y sky130_fd_sc_hd__a21oi_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2255_ hold865/X hold602/X _3466_/Q vssd1 vssd1 vccd1 vccd1 _2255_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2545__S1 _1942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2186_ _2661_/B _2200_/B vssd1 vssd1 vccd1 vccd1 _2201_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_79_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2870__A1 _2111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2075__B _2075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2790__S _2793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2030__S _2052_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3650__A _3659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2040_ _3507_/Q _3346_/Q vssd1 vssd1 vccd1 vccd1 _2040_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_76_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2942_ _3133_/A vssd1 vssd1 vccd1 vccd1 _2942_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2873_ hold594/X _2338_/B _2874_/S vssd1 vssd1 vccd1 vccd1 _2873_/X sky130_fd_sc_hd__mux2_1
X_1824_ _1824_/A _2383_/C vssd1 vssd1 vccd1 vccd1 _1831_/S sky130_fd_sc_hd__nand2_2
XFILLER_0_25_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1755_ _1811_/A _3566_/Q _1772_/B vssd1 vssd1 vccd1 vccd1 _1755_/X sky130_fd_sc_hd__or3_1
Xhold403 _2800_/X vssd1 vssd1 vccd1 vccd1 _3319_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold436 _3241_/Q vssd1 vssd1 vccd1 vccd1 hold436/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 _3300_/Q vssd1 vssd1 vccd1 vccd1 hold414/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 _2799_/X vssd1 vssd1 vccd1 vccd1 _3318_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 _2693_/X vssd1 vssd1 vccd1 vccd1 _3223_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 _2167_/X vssd1 vssd1 vccd1 vccd1 _3495_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold447 _3617_/Q vssd1 vssd1 vccd1 vccd1 _1571_/A sky130_fd_sc_hd__dlygate4sd3_1
X_1686_ hold100/X hold86/X hold21/X vssd1 vssd1 vccd1 vccd1 _3600_/D sky130_fd_sc_hd__mux2_1
X_3425_ _3427_/CLK _3425_/D vssd1 vssd1 vccd1 vccd1 _3425_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3356_ _3416_/CLK _3356_/D vssd1 vssd1 vccd1 vccd1 _3356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _3305_/CLK _3287_/D vssd1 vssd1 vccd1 vccd1 _3287_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2307_ hold357/X _2585_/A hold30/X vssd1 vssd1 vccd1 vccd1 _3444_/D sky130_fd_sc_hd__mux2_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2518__S1 _1911_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2238_ _2238_/A _2238_/B vssd1 vssd1 vccd1 vccd1 _2238_/Y sky130_fd_sc_hd__nor2_1
X_2169_ hold28/X _2410_/A _2169_/C vssd1 vssd1 vccd1 vccd1 _2661_/B sky130_fd_sc_hd__and3_4
XFILLER_0_63_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold970 _1764_/X vssd1 vssd1 vccd1 vccd1 _3563_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 _3345_/Q vssd1 vssd1 vccd1 vccd1 _2378_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold992 _3554_/Q vssd1 vssd1 vccd1 vccd1 _1744_/A sky130_fd_sc_hd__buf_1
XANTENNA__2785__S _2793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2770__A0 _2810_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3210_ _3331_/CLK _3210_/D vssd1 vssd1 vccd1 vccd1 _3210_/Q sky130_fd_sc_hd__dfxtp_1
X_3141_ _3612_/CLK _3141_/D vssd1 vssd1 vccd1 vccd1 _3141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3072_ _3073_/A vssd1 vssd1 vccd1 vccd1 _3072_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2825__A1 _2342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2023_ _2021_/X _2022_/X _2045_/S vssd1 vssd1 vccd1 vccd1 _2023_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_82_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2925_ _3095_/A vssd1 vssd1 vccd1 vccd1 _2925_/Y sky130_fd_sc_hd__inv_2
X_2856_ _2342_/B hold804/X _2864_/S vssd1 vssd1 vccd1 vccd1 _2856_/X sky130_fd_sc_hd__mux2_1
X_1807_ _1807_/A _1807_/B vssd1 vssd1 vccd1 vccd1 _3556_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2787_ _2807_/A1 hold214/X _2793_/S vssd1 vssd1 vccd1 vccd1 _2787_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold200 _1664_/X vssd1 vssd1 vccd1 vccd1 _3614_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 _2173_/Y vssd1 vssd1 vccd1 vccd1 _3494_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold233 _3316_/Q vssd1 vssd1 vccd1 vccd1 hold233/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 _2775_/X vssd1 vssd1 vccd1 vccd1 _3296_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1738_ _1851_/A _3456_/Q _1712_/Y _1718_/Y _1720_/Y vssd1 vssd1 vccd1 vccd1 _1741_/B
+ sky130_fd_sc_hd__o2111ai_1
Xhold244 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 input4/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 _2765_/X vssd1 vssd1 vccd1 vccd1 _3287_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 _2792_/X vssd1 vssd1 vccd1 vccd1 _3312_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 _3305_/Q vssd1 vssd1 vccd1 vccd1 hold255/X sky130_fd_sc_hd__dlygate4sd3_1
X_1669_ _1669_/A _2418_/B vssd1 vssd1 vccd1 vccd1 _2441_/A sky130_fd_sc_hd__nor2_2
Xhold299 _3445_/Q vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__dlygate4sd3_1
X_3408_ _3435_/CLK _3408_/D vssd1 vssd1 vccd1 vccd1 _3408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold288 _3616_/Q vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _3435_/CLK _3339_/D vssd1 vssd1 vccd1 vccd1 _3339_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2816__A1 _2097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2752__A0 _2812_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2807__A1 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2710_ _2810_/A1 hold315/X _2713_/S vssd1 vssd1 vccd1 vccd1 _2710_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2641_ _2824_/B _2905_/B _2875_/A vssd1 vssd1 vccd1 vccd1 _2650_/S sky130_fd_sc_hd__or3_4
XANTENNA__2743__A0 _2813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2572_ _2511_/Y _2581_/C _2571_/Y _2511_/B hold46/A vssd1 vssd1 vccd1 vccd1 _2573_/B
+ sky130_fd_sc_hd__a32o_1
XANTENNA__1607__B _1609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3124_ _3124_/A vssd1 vssd1 vccd1 vccd1 _3124_/Y sky130_fd_sc_hd__inv_2
X_3055_ _3055_/A vssd1 vssd1 vccd1 vccd1 _3055_/Y sky130_fd_sc_hd__inv_2
X_2006_ _1985_/S _2001_/X _2005_/X vssd1 vssd1 vccd1 vccd1 _2007_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__1769__S _3642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2908_ _2105_/A hold744/X _2914_/S vssd1 vssd1 vccd1 vccd1 _2908_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2839_ _2111_/B hold724/X _2843_/S vssd1 vssd1 vccd1 vccd1 _2839_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2725__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3493_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_output46_A _2580_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2624_ _2105_/B hold590/X _2629_/S vssd1 vssd1 vccd1 vccd1 _2624_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2716__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2555_ _2554_/X _2553_/X _3521_/Q vssd1 vssd1 vccd1 vccd1 _2556_/B sky130_fd_sc_hd__mux2_1
X_2486_ _2485_/X _2484_/X _2551_/S vssd1 vssd1 vccd1 vccd1 _2486_/X sky130_fd_sc_hd__mux2_1
X_3107_ _3114_/A vssd1 vssd1 vccd1 vccd1 _3107_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2168__B _3581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3038_ _3044_/A vssd1 vssd1 vccd1 vccd1 _3038_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_73_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2707__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold481_A _3581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2793__S _2793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput26 hold82/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__buf_1
XFILLER_0_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput37 input37/A vssd1 vssd1 vccd1 vccd1 _1907_/B sky130_fd_sc_hd__clkbuf_2
Xinput15 hold16/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3653__A _3659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2340_ _1569_/Y _2079_/A _2075_/B _1568_/Y vssd1 vssd1 vccd1 vccd1 _2344_/A sky130_fd_sc_hd__o22a_1
X_2271_ _2272_/B _2272_/C vssd1 vssd1 vccd1 vccd1 _2285_/B sky130_fd_sc_hd__and2_1
XANTENNA__2021__S1 _2044_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1986_ _3512_/Q _1985_/X _2052_/S vssd1 vssd1 vccd1 vccd1 _1986_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3656_ _3659_/A vssd1 vssd1 vccd1 vccd1 _3656_/X sky130_fd_sc_hd__buf_1
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout115_A _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2607_ _2338_/B hold766/X _2608_/S vssd1 vssd1 vccd1 vccd1 _2607_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3587_ _3614_/CLK _3587_/D _3078_/Y vssd1 vssd1 vccd1 vccd1 _3587_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2538_ hold70/A hold7/A vssd1 vssd1 vccd1 vccd1 _2538_/X sky130_fd_sc_hd__or2_1
X_2469_ _3370_/Q _3352_/Q _3361_/Q _3190_/Q _2554_/S0 _1911_/B vssd1 vssd1 vccd1 vccd1
+ _2469_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_78_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2788__S _2793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2003__S1 _2222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1840_ _1877_/A _1877_/B vssd1 vssd1 vccd1 vccd1 _1840_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_37_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1771_ _2111_/A vssd1 vssd1 vccd1 vccd1 _2381_/B sky130_fd_sc_hd__inv_2
X_3510_ _3513_/CLK _3510_/D _3004_/Y vssd1 vssd1 vccd1 vccd1 _3510_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold607 _2877_/X vssd1 vssd1 vccd1 vccd1 _3402_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 _3436_/Q vssd1 vssd1 vccd1 vccd1 hold618/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold629 _2608_/X vssd1 vssd1 vccd1 vccd1 _3151_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3441_ _3563_/CLK _3441_/D _2935_/Y vssd1 vssd1 vccd1 vccd1 _3441_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _3414_/CLK _3372_/D vssd1 vssd1 vccd1 vccd1 _3372_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _2323_/A _2323_/B vssd1 vssd1 vccd1 vccd1 _2323_/Y sky130_fd_sc_hd__xnor2_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2254_ hold843/X hold865/X _2258_/S vssd1 vssd1 vccd1 vccd1 _3472_/D sky130_fd_sc_hd__mux2_1
X_2185_ _2375_/B vssd1 vssd1 vccd1 vccd1 _2185_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_79_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1969_ hold353/X hold376/X hold327/X hold382/X _2224_/B _2193_/A1 vssd1 vssd1 vccd1
+ vccd1 _1969_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_55_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3639_ _3642_/CLK _3639_/D _3130_/Y vssd1 vssd1 vccd1 vccd1 _3639_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1992__S0 _1590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3637_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2377__A1 _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1983__S0 _2224_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold4 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2301__A1 hold52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2941_ _3133_/A vssd1 vssd1 vccd1 vccd1 _2941_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2872_ hold516/X _2075_/B _2874_/S vssd1 vssd1 vccd1 vccd1 _2872_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1823_ _1823_/A _1823_/B vssd1 vssd1 vccd1 vccd1 _3552_/D sky130_fd_sc_hd__nor2_1
XANTENNA__2368__A1 _2052_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1754_ _1751_/B _2383_/C _1753_/X vssd1 vssd1 vccd1 vccd1 _1754_/X sky130_fd_sc_hd__o21a_1
Xhold404 _3205_/Q vssd1 vssd1 vccd1 vccd1 hold404/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 _3239_/Q vssd1 vssd1 vccd1 vccd1 hold426/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold415 _2779_/X vssd1 vssd1 vccd1 vccd1 _3300_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 _3250_/Q vssd1 vssd1 vccd1 vccd1 hold459/X sky130_fd_sc_hd__dlygate4sd3_1
X_1685_ hold79/X hold33/X hold21/X vssd1 vssd1 vccd1 vccd1 _3601_/D sky130_fd_sc_hd__mux2_1
X_3424_ _3583_/CLK _3424_/D vssd1 vssd1 vccd1 vccd1 _3424_/Q sky130_fd_sc_hd__dfxtp_1
Xhold437 _2713_/X vssd1 vssd1 vccd1 vccd1 _3241_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold448 _3626_/Q vssd1 vssd1 vccd1 vccd1 _2054_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3355_ _3416_/CLK _3355_/D vssd1 vssd1 vccd1 vccd1 _3355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _3316_/CLK _3286_/D vssd1 vssd1 vccd1 vccd1 _3286_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ hold299/X _2395_/A hold30/X vssd1 vssd1 vccd1 vccd1 _3445_/D sky130_fd_sc_hd__mux2_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2237_ _3478_/Q _2241_/A _2260_/A vssd1 vssd1 vccd1 vccd1 _2237_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2168_ _3482_/Q _3581_/Q _2585_/B vssd1 vssd1 vccd1 vccd1 _2169_/C sky130_fd_sc_hd__and3b_1
XANTENNA__2891__S _2894_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2099_ _2062_/B _2088_/B _2089_/Y _2084_/B _2121_/A _1783_/A vssd1 vssd1 vccd1 vccd1
+ _2100_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_48_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout95_A _2193_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold960 _1899_/Y vssd1 vssd1 vccd1 vccd1 _3525_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 _3561_/Q vssd1 vssd1 vccd1 vccd1 hold971/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold982 _2372_/X vssd1 vssd1 vccd1 vccd1 _3345_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 _1819_/X vssd1 vssd1 vccd1 vccd1 _3554_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1970__S _2045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2522__B2 _2506_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2522__A1 _2583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3140_ _3513_/CLK _3140_/D vssd1 vssd1 vccd1 vccd1 _3140_/Q sky130_fd_sc_hd__dfxtp_1
X_3071_ _3073_/A vssd1 vssd1 vccd1 vccd1 _3071_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_82_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2022_ hold229/X hold257/X hold223/X hold248/X _2044_/S0 _2044_/S1 vssd1 vssd1 vccd1
+ vccd1 _2022_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2589__A1 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2924_ _3055_/A vssd1 vssd1 vccd1 vccd1 _2924_/Y sky130_fd_sc_hd__inv_2
X_2855_ _2885_/C _2875_/B vssd1 vssd1 vccd1 vccd1 _2864_/S sky130_fd_sc_hd__or2_4
XFILLER_0_72_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1806_ _1806_/A1 _1803_/B _1803_/A vssd1 vssd1 vccd1 vccd1 _1806_/Y sky130_fd_sc_hd__a21oi_1
X_2786_ _2806_/A1 hold187/X _2793_/S vssd1 vssd1 vccd1 vccd1 _2786_/X sky130_fd_sc_hd__mux2_1
Xhold201 _3599_/Q vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _2797_/X vssd1 vssd1 vccd1 vccd1 _3316_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1737_ _1881_/A _3446_/Q _1713_/Y _1714_/Y _1719_/Y vssd1 vssd1 vccd1 vccd1 _1741_/A
+ sky130_fd_sc_hd__o2111ai_1
XANTENNA__2761__A1 _2811_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold212 _3627_/Q vssd1 vssd1 vccd1 vccd1 _2081_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xhold223 _3199_/Q vssd1 vssd1 vccd1 vccd1 hold223/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 _3314_/Q vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 _2785_/X vssd1 vssd1 vccd1 vccd1 _3305_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 _3303_/Q vssd1 vssd1 vccd1 vccd1 hold278/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _1611_/X vssd1 vssd1 vccd1 vccd1 _1612_/B sky130_fd_sc_hd__dlygate4sd3_1
X_1668_ _1668_/A _2407_/A vssd1 vssd1 vccd1 vccd1 _2418_/B sky130_fd_sc_hd__nand2_1
XANTENNA__2886__S _2894_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3407_ _3523_/CLK _3407_/D vssd1 vssd1 vccd1 vccd1 _3407_/Q sky130_fd_sc_hd__dfxtp_1
Xhold289 _3613_/Q vssd1 vssd1 vccd1 vccd1 _1573_/A sky130_fd_sc_hd__dlygate4sd3_1
X_3338_ _3436_/CLK _3338_/D vssd1 vssd1 vccd1 vccd1 _3338_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1599_ _3346_/Q vssd1 vssd1 vccd1 vccd1 _2052_/S sky130_fd_sc_hd__clkinv_4
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3269_ _3305_/CLK _3269_/D vssd1 vssd1 vccd1 vccd1 _3269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold790 _3359_/Q vssd1 vssd1 vccd1 vccd1 hold790/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2097__A _2097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3656__A _3659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2640_ _2339_/B hold574/X _2640_/S vssd1 vssd1 vccd1 vccd1 _2640_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2571_ _2571_/A _2571_/B vssd1 vssd1 vccd1 vccd1 _2571_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3123_ _3126_/A vssd1 vssd1 vccd1 vccd1 _3123_/Y sky130_fd_sc_hd__inv_2
X_3054_ _3055_/A vssd1 vssd1 vccd1 vccd1 _3054_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2005_ _1985_/S _2005_/B vssd1 vssd1 vccd1 vccd1 _2005_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2907_ _2097_/A hold742/X _2914_/S vssd1 vssd1 vccd1 vccd1 _2907_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2838_ _2105_/B hold698/X _2843_/S vssd1 vssd1 vccd1 vccd1 _2838_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2769_ _2809_/A1 hold388/X _2773_/S vssd1 vssd1 vccd1 vccd1 _2769_/X sky130_fd_sc_hd__mux2_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2670__A0 _2811_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output39_A _3443_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2623_ _2105_/A hold682/X _2629_/S vssd1 vssd1 vccd1 vccd1 _2623_/X sky130_fd_sc_hd__mux2_1
X_2554_ _3178_/Q _3427_/Q _3418_/Q _3160_/Q _2554_/S0 _1942_/A vssd1 vssd1 vccd1 vccd1
+ _2554_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_50_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2485_ _3182_/Q _3335_/Q _3164_/Q _3146_/Q _1943_/B _2550_/S1 vssd1 vssd1 vccd1 vccd1
+ _2485_/X sky130_fd_sc_hd__mux4_1
X_3106_ _3114_/A vssd1 vssd1 vccd1 vccd1 _3106_/Y sky130_fd_sc_hd__inv_2
X_3037_ _3044_/A vssd1 vssd1 vccd1 vccd1 _3037_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2652__A0 _2342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_46_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3414_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2643__A0 _2097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput27 input27/A vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_2
Xinput16 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 _1625_/B sky130_fd_sc_hd__buf_2
XFILLER_0_12_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2270_ _1889_/Y _2269_/X _2272_/C vssd1 vssd1 vccd1 vccd1 _2285_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_74_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1685__A1 hold33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2882__A0 _2075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2634__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1985_ _1984_/X _1981_/X _1985_/S vssd1 vssd1 vccd1 vccd1 _1985_/X sky130_fd_sc_hd__mux2_2
X_3655_ _3659_/A vssd1 vssd1 vccd1 vccd1 _3655_/X sky130_fd_sc_hd__buf_1
XFILLER_0_2_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2606_ _2075_/B hold588/X _2608_/S vssd1 vssd1 vccd1 vccd1 _2606_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout108_A hold123/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3586_ _3609_/CLK _3586_/D _3077_/Y vssd1 vssd1 vccd1 vccd1 _3586_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2537_ hold68/A _2568_/B _2417_/B _3379_/Q _2536_/X vssd1 vssd1 vccd1 vccd1 _2537_/X
+ sky130_fd_sc_hd__o221a_1
X_2468_ _2467_/X _2466_/X _2551_/S vssd1 vssd1 vccd1 vccd1 _2468_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2894__S _2894_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2399_ hold33/X _2403_/B vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__and2_1
XANTENNA__2625__A0 _2111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1973__S _2045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2864__A0 _2339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1667__A1 _2585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2616__A0 _2075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2552__B _3522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1770_ _1769_/X _3443_/Q _1770_/S vssd1 vssd1 vccd1 vccd1 _2111_/A sky130_fd_sc_hd__mux2_4
XFILLER_0_64_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold608 _3170_/Q vssd1 vssd1 vccd1 vccd1 hold608/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold619 _2914_/X vssd1 vssd1 vccd1 vccd1 _3436_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3440_ _3563_/CLK _3440_/D _2934_/Y vssd1 vssd1 vccd1 vccd1 _3440_/Q sky130_fd_sc_hd__dfrtp_1
X_3371_ _3423_/CLK _3371_/D vssd1 vssd1 vccd1 vccd1 _3371_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2322_ _2322_/A _2322_/B vssd1 vssd1 vccd1 vccd1 _2323_/B sky130_fd_sc_hd__xnor2_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2253_ hold812/X hold843/X _3466_/Q vssd1 vssd1 vccd1 vccd1 _2253_/X sky130_fd_sc_hd__mux2_1
X_2184_ _2145_/A _2183_/X _2366_/B _2366_/A vssd1 vssd1 vccd1 vccd1 _2200_/B sky130_fd_sc_hd__o211ai_4
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__2607__A0 _2338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1968_ hold408/X hold345/X hold396/X hold341/X _2044_/S0 _2044_/S1 vssd1 vssd1 vccd1
+ vccd1 _1968_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_55_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2889__S _2894_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1899_ _1897_/X _1898_/Y _1933_/A vssd1 vssd1 vccd1 vccd1 _1899_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3638_ _3642_/CLK _3638_/D _3129_/Y vssd1 vssd1 vccd1 vccd1 _3638_/Q sky130_fd_sc_hd__dfrtp_1
X_3569_ _3571_/CLK _3569_/D _3063_/Y vssd1 vssd1 vccd1 vccd1 _3569_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__1992__S1 _2222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2846__A0 _2097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1649__A1 hold44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1983__S1 _2222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2837__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__buf_1
XANTENNA__3659__A _3659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2940_ _3128_/A vssd1 vssd1 vccd1 vccd1 _2940_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_84_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2871_ hold556/X _2079_/A _2874_/S vssd1 vssd1 vccd1 vccd1 _2871_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1822_ _1810_/A _1817_/B _1817_/A vssd1 vssd1 vccd1 vccd1 _1823_/B sky130_fd_sc_hd__o21a_1
X_1753_ _1811_/A _3567_/Q _1772_/B vssd1 vssd1 vccd1 vccd1 _1753_/X sky130_fd_sc_hd__or3_1
XFILLER_0_80_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1684_ hold78/X hold52/X hold21/X vssd1 vssd1 vccd1 vccd1 _3602_/D sky130_fd_sc_hd__mux2_1
Xhold405 _2672_/X vssd1 vssd1 vccd1 vccd1 _3205_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 _2711_/X vssd1 vssd1 vccd1 vccd1 _3239_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 _3257_/Q vssd1 vssd1 vccd1 vccd1 hold416/X sky130_fd_sc_hd__dlygate4sd3_1
X_3423_ _3423_/CLK _3423_/D vssd1 vssd1 vccd1 vccd1 _3423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold449 _1642_/X vssd1 vssd1 vccd1 vccd1 _3626_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 _3309_/Q vssd1 vssd1 vccd1 vccd1 hold438/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _3414_/CLK _3354_/D vssd1 vssd1 vccd1 vccd1 _3354_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ hold444/X _2396_/A hold30/X vssd1 vssd1 vccd1 vccd1 _3446_/D sky130_fd_sc_hd__mux2_1
X_3285_ _3316_/CLK _3285_/D vssd1 vssd1 vccd1 vccd1 _3285_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2236_ _2236_/A _2236_/B vssd1 vssd1 vccd1 vccd1 _2236_/X sky130_fd_sc_hd__and2_1
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2167_ _3495_/Q _1931_/B _2166_/Y _1933_/A vssd1 vssd1 vccd1 vccd1 _2167_/X sky130_fd_sc_hd__a211o_1
X_2098_ _2339_/B _2098_/B vssd1 vssd1 vccd1 vccd1 _2106_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold972 _1768_/X vssd1 vssd1 vccd1 vccd1 _3561_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 _3501_/Q vssd1 vssd1 vccd1 vccd1 _2134_/B sky130_fd_sc_hd__clkbuf_2
Xhold950 _1752_/X vssd1 vssd1 vccd1 vccd1 _3569_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout88_A _1911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold994 _3555_/Q vssd1 vssd1 vccd1 vccd1 _1745_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold983 _3570_/Q vssd1 vssd1 vccd1 vccd1 hold983/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3070_ _3070_/A vssd1 vssd1 vccd1 vccd1 _3070_/Y sky130_fd_sc_hd__inv_2
X_2021_ hold272/X hold274/X hold227/X hold235/X _2044_/S0 _2044_/S1 vssd1 vssd1 vccd1
+ vccd1 _2021_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_82_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2923_ _3133_/A vssd1 vssd1 vccd1 vccd1 _2923_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2854_ _3526_/Q _2905_/B vssd1 vssd1 vccd1 vccd1 _2875_/B sky130_fd_sc_hd__nand2_2
X_2785_ _2805_/A1 hold255/X _2793_/S vssd1 vssd1 vccd1 vccd1 _2785_/X sky130_fd_sc_hd__mux2_1
X_1805_ _1803_/B _1804_/X _1807_/A _1797_/B vssd1 vssd1 vccd1 vccd1 _3557_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_31_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1736_ _1743_/B _1743_/C vssd1 vssd1 vccd1 vccd1 _2231_/B sky130_fd_sc_hd__nor2_1
Xhold202 _3135_/Q vssd1 vssd1 vccd1 vccd1 hold202/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 _1641_/X vssd1 vssd1 vccd1 vccd1 _3627_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 _3226_/Q vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _2666_/X vssd1 vssd1 vccd1 vccd1 _3199_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 _2795_/X vssd1 vssd1 vccd1 vccd1 _3314_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1667_ _1575_/A _2585_/A _1667_/S vssd1 vssd1 vccd1 vccd1 _3611_/D sky130_fd_sc_hd__mux2_1
Xhold257 _3208_/Q vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 _2661_/B vssd1 vssd1 vccd1 vccd1 _2587_/C sky130_fd_sc_hd__buf_2
Xhold279 _2782_/X vssd1 vssd1 vccd1 vccd1 _3303_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3406_ _3435_/CLK _3406_/D vssd1 vssd1 vccd1 vccd1 _3406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1598_ _3341_/Q vssd1 vssd1 vccd1 vccd1 _1598_/Y sky130_fd_sc_hd__inv_2
X_3337_ _3435_/CLK _3337_/D vssd1 vssd1 vccd1 vccd1 _3337_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _3316_/CLK _3268_/D vssd1 vssd1 vccd1 vccd1 _3268_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2219_ _2207_/B _2214_/Y _2218_/X _2214_/B _2205_/A vssd1 vssd1 vccd1 vccd1 _2219_/X
+ sky130_fd_sc_hd__a32o_1
X_3199_ _3325_/CLK _3199_/D vssd1 vssd1 vccd1 vccd1 _3199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1981__S _2045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold780 _3166_/Q vssd1 vssd1 vccd1 vccd1 hold780/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 _2835_/X vssd1 vssd1 vccd1 vccd1 _3359_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2097__B _2342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2052__S _2052_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2570_ _2583_/B _2570_/B vssd1 vssd1 vccd1 vccd1 _2570_/X sky130_fd_sc_hd__and2_2
XFILLER_0_50_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3122_ _3133_/A vssd1 vssd1 vccd1 vccd1 _3122_/Y sky130_fd_sc_hd__inv_2
X_3053_ _3055_/A vssd1 vssd1 vccd1 vccd1 _3053_/Y sky130_fd_sc_hd__inv_2
X_2004_ _2003_/X _2002_/X _2045_/S vssd1 vssd1 vccd1 vccd1 _2005_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2906_ _2342_/B hold558/X _2914_/S vssd1 vssd1 vccd1 vccd1 _2906_/X sky130_fd_sc_hd__mux2_1
X_2837_ _2105_/A hold700/X _2843_/S vssd1 vssd1 vccd1 vccd1 _2837_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2768_ _2808_/A1 hold157/X _2773_/S vssd1 vssd1 vccd1 vccd1 _2768_/X sky130_fd_sc_hd__mux2_1
X_1719_ _3541_/Q _3458_/Q vssd1 vssd1 vccd1 vccd1 _1719_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__2897__S _2904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2699_ _2809_/A1 hold400/X _2703_/S vssd1 vssd1 vccd1 vccd1 _2699_/X sky130_fd_sc_hd__mux2_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2033__S0 _2044_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2622_ _2097_/A hold632/X _2629_/S vssd1 vssd1 vccd1 vccd1 _2622_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2553_ _3376_/Q _3358_/Q _3367_/Q _3196_/Q _2554_/S0 _1911_/B vssd1 vssd1 vccd1 vccd1
+ _2553_/X sky130_fd_sc_hd__mux4_1
X_2484_ _3404_/Q _3395_/Q _3386_/Q _3431_/Q _1943_/B _2550_/S1 vssd1 vssd1 vccd1 vccd1
+ _2484_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2024__S0 _1590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3105_ _3105_/A vssd1 vssd1 vccd1 vccd1 _3105_/Y sky130_fd_sc_hd__inv_2
X_3036_ _3036_/A vssd1 vssd1 vccd1 vccd1 _3036_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3483_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout70_A _2109_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2340__B1 _2075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput17 hold64/X vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__buf_2
Xinput28 input28/A vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_1
XFILLER_0_24_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2566__A _2583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2505__S _3522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1984_ _1983_/X _1982_/X _2045_/S vssd1 vssd1 vccd1 vccd1 _1984_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3654_ _3659_/A vssd1 vssd1 vccd1 vccd1 _3654_/X sky130_fd_sc_hd__buf_1
XFILLER_0_15_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2605_ _2079_/A hold754/X _2608_/S vssd1 vssd1 vccd1 vccd1 _2605_/X sky130_fd_sc_hd__mux2_1
X_3585_ _3633_/CLK _3585_/D _3076_/Y vssd1 vssd1 vccd1 vccd1 _3585_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2536_ _3591_/Q hold67/A vssd1 vssd1 vccd1 vccd1 _2536_/X sky130_fd_sc_hd__or2_1
X_2467_ _3181_/Q _3334_/Q _3163_/Q _3145_/Q _1943_/B _2550_/S1 vssd1 vssd1 vccd1 vccd1
+ _2467_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2398_ hold86/X _2403_/B vssd1 vssd1 vccd1 vccd1 _3588_/D sky130_fd_sc_hd__and2_1
XFILLER_0_3_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2873__A1 _2338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3019_ _3089_/A vssd1 vssd1 vccd1 vccd1 _3019_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_38_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3100__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2484__S0 _1943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2561__B1 _2506_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold609 _2632_/X vssd1 vssd1 vccd1 vccd1 _3170_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3370_ _3582_/CLK _3370_/D vssd1 vssd1 vccd1 vccd1 _3370_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2321_ _1966_/B _2321_/B vssd1 vssd1 vccd1 vccd1 _2322_/B sky130_fd_sc_hd__and2b_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2252_ _2252_/A0 hold812/X _3466_/Q vssd1 vssd1 vccd1 vccd1 _2252_/X sky130_fd_sc_hd__mux2_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2183_ _2383_/A _3345_/Q vssd1 vssd1 vccd1 vccd1 _2183_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_26_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2466__S0 _1943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1967_ hold822/X _1966_/Y _2053_/S vssd1 vssd1 vccd1 vccd1 _1967_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout120_A _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2791__A0 _2811_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1898_ _2905_/B _2630_/C vssd1 vssd1 vccd1 vccd1 _1898_/Y sky130_fd_sc_hd__nand2_1
X_3637_ _3637_/CLK hold39/X _3128_/Y vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3568_ _3571_/CLK _3568_/D _3062_/Y vssd1 vssd1 vccd1 vccd1 _3568_/Q sky130_fd_sc_hd__dfstp_1
X_2519_ _3175_/Q _3424_/Q _3415_/Q _3157_/Q _2554_/S0 _1911_/B vssd1 vssd1 vccd1 vccd1
+ _2519_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3499_ _3499_/CLK _3499_/D _2993_/Y vssd1 vssd1 vccd1 vccd1 _3499_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_66_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1984__S _2045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2782__A0 _2812_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3631_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2870_ hold680/X _2111_/B _2874_/S vssd1 vssd1 vccd1 vccd1 _2870_/X sky130_fd_sc_hd__mux2_1
X_1821_ _1774_/C _1823_/A _1821_/B1 _1817_/B vssd1 vssd1 vccd1 vccd1 _1821_/X sky130_fd_sc_hd__o22a_1
XANTENNA__2448__S0 _1943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2773__A0 _2813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1752_ _1749_/B _2383_/C _1751_/X vssd1 vssd1 vccd1 vccd1 _1752_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_40_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1907__B _1907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold417 _2731_/X vssd1 vssd1 vccd1 vccd1 _3257_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold406 _3138_/Q vssd1 vssd1 vccd1 vccd1 hold406/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1683_ hold68/X hold44/X hold21/X vssd1 vssd1 vccd1 vccd1 _3603_/D sky130_fd_sc_hd__mux2_1
X_3422_ _3423_/CLK _3422_/D vssd1 vssd1 vccd1 vccd1 _3422_/Q sky130_fd_sc_hd__dfxtp_1
Xhold428 _3210_/Q vssd1 vssd1 vccd1 vccd1 hold428/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 _2789_/X vssd1 vssd1 vccd1 vccd1 _3309_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _3423_/CLK _3353_/D vssd1 vssd1 vccd1 vccd1 _3353_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _3319_/CLK _3284_/D vssd1 vssd1 vccd1 vccd1 _3284_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ hold204/X _2397_/A hold30/X vssd1 vssd1 vccd1 vccd1 _3447_/D sky130_fd_sc_hd__mux2_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2828__A1 _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2235_ _2261_/A _2238_/A _2261_/B vssd1 vssd1 vccd1 vccd1 _2235_/X sky130_fd_sc_hd__a21o_1
X_2166_ _2162_/X _2163_/Y _2165_/X _1922_/B _2598_/C vssd1 vssd1 vccd1 vccd1 _2166_/Y
+ sky130_fd_sc_hd__a2111oi_1
X_2097_ _2097_/A _2342_/B vssd1 vssd1 vccd1 vccd1 _2098_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2999_ _3121_/A vssd1 vssd1 vccd1 vccd1 _2999_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold940 _3504_/Q vssd1 vssd1 vccd1 vccd1 _1588_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold962 _2140_/Y vssd1 vssd1 vccd1 vccd1 hold962/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 _3566_/Q vssd1 vssd1 vccd1 vccd1 hold973/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold951 _3498_/Q vssd1 vssd1 vccd1 vccd1 _2130_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 _1816_/X vssd1 vssd1 vccd1 vccd1 _3555_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 _1750_/X vssd1 vssd1 vccd1 vccd1 _3570_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2819__A1 _2111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2020_ hold814/X _2019_/Y _2053_/S vssd1 vssd1 vccd1 vccd1 _2020_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_82_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2922_ _3065_/A vssd1 vssd1 vccd1 vccd1 _2922_/Y sky130_fd_sc_hd__inv_2
X_2853_ _2339_/B hold634/X _2853_/S vssd1 vssd1 vccd1 vccd1 _2853_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1804_ _1797_/B _1803_/A _1604_/Y vssd1 vssd1 vccd1 vccd1 _1804_/X sky130_fd_sc_hd__a21o_1
X_2784_ _2794_/A _2794_/B _2784_/C vssd1 vssd1 vccd1 vccd1 _2793_/S sky130_fd_sc_hd__or3_4
XANTENNA__2746__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1735_ _1735_/A _1735_/B _1735_/C _1735_/D vssd1 vssd1 vccd1 vccd1 _1743_/C sky130_fd_sc_hd__or4_2
XFILLER_0_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold214 _3307_/Q vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 _3242_/Q vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 _2590_/X vssd1 vssd1 vccd1 vccd1 _3135_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 _3276_/Q vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1666_ _1574_/A _2395_/A _1667_/S vssd1 vssd1 vccd1 vccd1 _3612_/D sky130_fd_sc_hd__mux2_1
Xhold258 _2676_/X vssd1 vssd1 vccd1 vccd1 _3208_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 _2697_/X vssd1 vssd1 vccd1 vccd1 _3226_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 _2182_/X vssd1 vssd1 vccd1 vccd1 _3491_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1597_ _3342_/Q vssd1 vssd1 vccd1 vccd1 _1597_/Y sky130_fd_sc_hd__inv_2
X_3405_ _3435_/CLK _3405_/D vssd1 vssd1 vccd1 vccd1 _3405_/Q sky130_fd_sc_hd__dfxtp_1
X_3336_ _3404_/CLK _3336_/D vssd1 vssd1 vccd1 vccd1 _3336_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _3316_/CLK _3267_/D vssd1 vssd1 vccd1 vccd1 _3267_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2218_ _3483_/Q _2218_/B vssd1 vssd1 vccd1 vccd1 _2218_/X sky130_fd_sc_hd__or2_1
X_3198_ _3328_/CLK _3198_/D vssd1 vssd1 vccd1 vccd1 _3198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2149_ _2149_/A _2149_/B vssd1 vssd1 vccd1 vccd1 _2149_/X sky130_fd_sc_hd__or2_1
XANTENNA__2737__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold781 _2626_/X vssd1 vssd1 vccd1 vccd1 _3166_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold770 _3354_/Q vssd1 vssd1 vccd1 vccd1 hold770/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 _3184_/Q vssd1 vssd1 vccd1 vccd1 hold792/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2394__A _2585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2728__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3121_ _3121_/A vssd1 vssd1 vccd1 vccd1 _3121_/Y sky130_fd_sc_hd__inv_2
X_3052_ _3070_/A vssd1 vssd1 vccd1 vccd1 _3052_/Y sky130_fd_sc_hd__inv_2
X_2003_ hold420/X _3318_/Q hold438/X hold414/X _2224_/B _2222_/A vssd1 vssd1 vccd1
+ vccd1 _2003_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_77_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2905_ _3526_/Q _2905_/B _2905_/C vssd1 vssd1 vccd1 vccd1 _2914_/S sky130_fd_sc_hd__nand3_4
X_2836_ _2097_/A hold702/X _2843_/S vssd1 vssd1 vccd1 vccd1 _2836_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2719__A0 _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2767_ _2807_/A1 hold219/X _2773_/S vssd1 vssd1 vccd1 vccd1 _2767_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1718_ _3445_/Q _1883_/A vssd1 vssd1 vccd1 vccd1 _1718_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_13_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2698_ _2808_/A1 hold138/X _2703_/S vssd1 vssd1 vccd1 vccd1 _2698_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1649_ hold69/X hold44/X hold60/X vssd1 vssd1 vccd1 vccd1 _3622_/D sky130_fd_sc_hd__mux2_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ _3319_/CLK _3319_/D vssd1 vssd1 vccd1 vccd1 _3319_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2033__S1 _2044_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2343__D1 _1889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2621_ _2342_/B hold774/X _2629_/S vssd1 vssd1 vccd1 vccd1 _2621_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2552_ _2551_/X _3522_/Q vssd1 vssd1 vccd1 vccd1 _2552_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_10_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2483_ _3447_/Q hold29/A _2583_/B _2482_/X vssd1 vssd1 vccd1 vccd1 _2483_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2024__S1 _2222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3104_ _3105_/A vssd1 vssd1 vccd1 vccd1 _3104_/Y sky130_fd_sc_hd__inv_2
X_3035_ _3036_/A vssd1 vssd1 vccd1 vccd1 _3035_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2819_ hold536/X _2111_/B _2823_/S vssd1 vssd1 vccd1 vccd1 _2819_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1987__S _2053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput18 input18/A vssd1 vssd1 vccd1 vccd1 _1660_/A sky130_fd_sc_hd__clkbuf_2
Xinput29 input29/A vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_1
XANTENNA__2611__S _2618_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output44_A _2576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1983_ _3248_/Q _3320_/Q _3311_/Q _3302_/Q _2224_/B _2222_/A vssd1 vssd1 vccd1 vccd1
+ _1983_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3653_ _3659_/A vssd1 vssd1 vccd1 vccd1 _3653_/X sky130_fd_sc_hd__buf_1
XANTENNA__2521__S _3522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2604_ _2111_/B hold738/X _2608_/S vssd1 vssd1 vccd1 vccd1 _2604_/X sky130_fd_sc_hd__mux2_1
X_3584_ _3609_/CLK _3584_/D _3075_/Y vssd1 vssd1 vccd1 vccd1 _3584_/Q sky130_fd_sc_hd__dfrtp_1
X_2535_ _2583_/B _2527_/X _2534_/X _2506_/S vssd1 vssd1 vccd1 vccd1 _2535_/X sky130_fd_sc_hd__a22o_1
X_2466_ _3403_/Q _3394_/Q _3385_/Q _3430_/Q _1943_/B _2550_/S1 vssd1 vssd1 vccd1 vccd1
+ _2466_/X sky130_fd_sc_hd__mux4_1
X_2397_ _2397_/A _2403_/B vssd1 vssd1 vccd1 vccd1 _3587_/D sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3018_ _3089_/A vssd1 vssd1 vccd1 vccd1 _3018_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_58_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2484__S1 _2550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1994__A_N _1985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2561__A1 _1595_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2320_ _2318_/X _2319_/X _2320_/S vssd1 vssd1 vccd1 vccd1 _2322_/A sky130_fd_sc_hd__mux2_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2251_ hold602/X _2248_/X _2250_/X _3475_/Q vssd1 vssd1 vccd1 vccd1 _2251_/X sky130_fd_sc_hd__a22o_1
XANTENNA__2304__A1 _2397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2182_ _3491_/Q _2587_/C _2181_/Y vssd1 vssd1 vccd1 vccd1 _2182_/X sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_0_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3433_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1966_ _3346_/Q _1966_/B vssd1 vssd1 vccd1 vccd1 _1966_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2466__S1 _2550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1897_ _2630_/C _1945_/B _1945_/C vssd1 vssd1 vccd1 vccd1 _1897_/X sky130_fd_sc_hd__or3_1
X_3636_ _3636_/CLK _3636_/D _3127_/Y vssd1 vssd1 vccd1 vccd1 _3636_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout113_A hold176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3567_ _3580_/CLK _3567_/D _3061_/Y vssd1 vssd1 vccd1 vccd1 _3567_/Q sky130_fd_sc_hd__dfstp_1
X_2518_ _3373_/Q _3355_/Q _3364_/Q _3193_/Q _2554_/S0 _1911_/B vssd1 vssd1 vccd1 vccd1
+ _2518_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_11_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3498_ _3499_/CLK _3498_/D _2992_/Y vssd1 vssd1 vccd1 vccd1 _3498_/Q sky130_fd_sc_hd__dfrtp_1
X_2449_ _3180_/Q _3333_/Q _3162_/Q _3144_/Q _1943_/B _2550_/S1 vssd1 vssd1 vccd1 vccd1
+ _2449_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1968__S0 _2044_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2397__A _2397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1820_ _1774_/C _1580_/A _1810_/A vssd1 vssd1 vccd1 vccd1 _1820_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__2448__S1 _1942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1751_ _1811_/A _1751_/B _1772_/B vssd1 vssd1 vccd1 vccd1 _1751_/X sky130_fd_sc_hd__or3_1
Xhold418 _3331_/Q vssd1 vssd1 vccd1 vccd1 hold418/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold407 _2593_/X vssd1 vssd1 vccd1 vccd1 _3138_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1682_ hold74/X hold49/X hold21/X vssd1 vssd1 vccd1 vccd1 _3604_/D sky130_fd_sc_hd__mux2_1
X_3421_ _3583_/CLK _3421_/D vssd1 vssd1 vccd1 vccd1 _3421_/Q sky130_fd_sc_hd__dfxtp_1
Xhold429 _2678_/X vssd1 vssd1 vccd1 vccd1 _3210_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3352_ _3369_/CLK _3352_/D vssd1 vssd1 vccd1 vccd1 _3352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1959__S0 _2044_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ hold88/X hold86/X hold30/X vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__mux2_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _3305_/CLK _3283_/D vssd1 vssd1 vccd1 vccd1 _3283_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ _2261_/A _2236_/A vssd1 vssd1 vccd1 vccd1 _2234_/Y sky130_fd_sc_hd__xnor2_1
X_2165_ _2165_/A _2165_/B _1944_/B vssd1 vssd1 vccd1 vccd1 _2165_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_45_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2096_ _2059_/A _2080_/B _2095_/X _2067_/B vssd1 vssd1 vccd1 vccd1 _2096_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_0_48_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2998_ _3121_/A vssd1 vssd1 vccd1 vccd1 _2998_/Y sky130_fd_sc_hd__inv_2
X_1949_ _1891_/A _1948_/Y _1910_/B vssd1 vssd1 vccd1 vccd1 _1949_/X sky130_fd_sc_hd__o21a_1
Xhold930 _2385_/X vssd1 vssd1 vccd1 vccd1 _3440_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3619_ _3631_/CLK _3619_/D _3110_/Y vssd1 vssd1 vccd1 vccd1 _3619_/Q sky130_fd_sc_hd__dfrtp_1
Xhold963 _2142_/Y vssd1 vssd1 vccd1 vccd1 _3501_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 _2120_/Y vssd1 vssd1 vccd1 vccd1 _3504_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold952 _2155_/X vssd1 vssd1 vccd1 vccd1 hold952/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 _3533_/Q vssd1 vssd1 vccd1 vccd1 _1843_/A sky130_fd_sc_hd__buf_1
Xhold996 _3541_/Q vssd1 vssd1 vccd1 vccd1 _1853_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold974 _1758_/X vssd1 vssd1 vccd1 vccd1 _3566_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2755__A1 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2691__A0 _2811_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2921_ _3065_/A vssd1 vssd1 vccd1 vccd1 _2921_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2852_ _2338_/B hold778/X _2853_/S vssd1 vssd1 vccd1 vccd1 _2852_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2783_ _2813_/A1 hold378/X _2783_/S vssd1 vssd1 vccd1 vccd1 _2783_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1803_ _1803_/A _1803_/B vssd1 vssd1 vccd1 vccd1 _1807_/A sky130_fd_sc_hd__and2_1
X_1734_ _1871_/A _1596_/Y hold444/X _1881_/A _1725_/X vssd1 vssd1 vccd1 vccd1 _1735_/D
+ sky130_fd_sc_hd__a221o_1
Xhold215 _2787_/X vssd1 vssd1 vccd1 vccd1 _3307_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 _2715_/X vssd1 vssd1 vccd1 vccd1 _3242_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 _3447_/Q vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 _3271_/Q vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
X_3404_ _3404_/CLK _3404_/D vssd1 vssd1 vccd1 vccd1 _3404_/Q sky130_fd_sc_hd__dfxtp_1
X_1665_ _1573_/A _2396_/A _1667_/S vssd1 vssd1 vccd1 vccd1 _3613_/D sky130_fd_sc_hd__mux2_1
Xhold259 _3493_/Q vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 _3325_/Q vssd1 vssd1 vccd1 vccd1 hold248/X sky130_fd_sc_hd__dlygate4sd3_1
X_1596_ hold62/X vssd1 vssd1 vccd1 vccd1 _1596_/Y sky130_fd_sc_hd__inv_2
X_3335_ _3404_/CLK _3335_/D vssd1 vssd1 vccd1 vccd1 _3335_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ _3488_/CLK _3266_/D vssd1 vssd1 vccd1 vccd1 _3266_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2217_ _2212_/B _2214_/Y _2216_/X _2214_/B _2208_/A vssd1 vssd1 vccd1 vccd1 _2217_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2187__D _2200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3197_ _3325_/CLK _3197_/D vssd1 vssd1 vccd1 vccd1 _3197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2148_ _2149_/A _2149_/B vssd1 vssd1 vccd1 vccd1 _2156_/B sky130_fd_sc_hd__nor2_2
X_2079_ _2079_/A _2079_/B vssd1 vssd1 vccd1 vccd1 _2107_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold782 _3406_/Q vssd1 vssd1 vccd1 vccd1 hold782/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 _2829_/X vssd1 vssd1 vccd1 vccd1 _3354_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold760 _3154_/Q vssd1 vssd1 vccd1 vccd1 hold760/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold793 _2647_/X vssd1 vssd1 vccd1 vccd1 _3184_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2614__S _2618_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2900__A1 _2109_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3120_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3120_/Y sky130_fd_sc_hd__inv_2
X_3051_ _3070_/A vssd1 vssd1 vccd1 vccd1 _3051_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2585__A _2585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2002_ _3291_/Q _3282_/Q _3273_/Q _3264_/Q _2044_/S0 _2044_/S1 vssd1 vssd1 vccd1
+ vccd1 _2002_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2664__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2904_ hold530/X _2081_/X _2904_/S vssd1 vssd1 vccd1 vccd1 _2904_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2835_ _2342_/B hold790/X _2843_/S vssd1 vssd1 vccd1 vccd1 _2835_/X sky130_fd_sc_hd__mux2_1
X_2766_ _2806_/A1 hold167/X _2773_/S vssd1 vssd1 vccd1 vccd1 _2766_/X sky130_fd_sc_hd__mux2_1
X_1717_ hold88/A _3531_/Q vssd1 vssd1 vccd1 vccd1 _1717_/X sky130_fd_sc_hd__and2b_1
X_2697_ _2807_/A1 hold235/X _2703_/S vssd1 vssd1 vccd1 vccd1 _2697_/X sky130_fd_sc_hd__mux2_1
X_1648_ _3623_/Q hold49/X hold60/A vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__mux2_1
XFILLER_0_6_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1579_ _3607_/Q vssd1 vssd1 vccd1 vccd1 _1579_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3318_ _3318_/CLK _3318_/D vssd1 vssd1 vccd1 vccd1 _3318_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3249_ _3488_/CLK _3249_/D vssd1 vssd1 vccd1 vccd1 _3249_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2655__A0 _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2502__S0 _1943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2434__S _3522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold590 _3164_/Q vssd1 vssd1 vccd1 vccd1 hold590/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2646__A0 _2111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1621__A1 _2396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2620_ _2824_/B _2905_/B _2885_/C vssd1 vssd1 vccd1 vccd1 _2629_/S sky130_fd_sc_hd__or3_4
XFILLER_0_2_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2551_ _2550_/X _2549_/X _2551_/S vssd1 vssd1 vccd1 vccd1 _2551_/X sky130_fd_sc_hd__mux2_1
X_2482_ _3641_/Q _2511_/A _2511_/B _2481_/X vssd1 vssd1 vccd1 vccd1 _2482_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_50_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1688__A1 _2396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold14_A hold14/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3103_ _3105_/A vssd1 vssd1 vccd1 vccd1 _3103_/Y sky130_fd_sc_hd__inv_2
X_3034_ _3036_/A vssd1 vssd1 vccd1 vccd1 _3034_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2637__A0 _2079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1659__A _1659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2818_ hold550/X _2105_/B _2823_/S vssd1 vssd1 vccd1 vccd1 _2818_/X sky130_fd_sc_hd__mux2_1
X_2749_ _2809_/A1 hold339/X _2753_/S vssd1 vssd1 vccd1 vccd1 _2749_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2876__A0 _2342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2340__A2 _2079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2628__A0 _2338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3539_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xinput19 input19/A vssd1 vssd1 vccd1 vccd1 _1609_/B sky130_fd_sc_hd__buf_2
XFILLER_0_20_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1982_ _3293_/Q _3284_/Q _3275_/Q _3266_/Q _1590_/A _2193_/A1 vssd1 vssd1 vccd1 vccd1
+ _1982_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_7_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3652_ _3659_/A vssd1 vssd1 vccd1 vccd1 _3652_/X sky130_fd_sc_hd__buf_1
X_2603_ _2105_/B hold716/X _2608_/S vssd1 vssd1 vccd1 vccd1 _2603_/X sky130_fd_sc_hd__mux2_1
X_3583_ _3583_/CLK _3583_/D vssd1 vssd1 vccd1 vccd1 _3583_/Q sky130_fd_sc_hd__dfxtp_1
X_2534_ _2533_/X _2530_/X _3522_/Q vssd1 vssd1 vccd1 vccd1 _2534_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1942__A _1942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2465_ _3446_/Q hold29/A _2456_/X _2464_/X _2583_/B vssd1 vssd1 vccd1 vccd1 _2465_/X
+ sky130_fd_sc_hd__o221a_1
X_2396_ _2396_/A _2403_/B vssd1 vssd1 vccd1 vccd1 _2396_/X sky130_fd_sc_hd__and2_1
XANTENNA__2858__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3017_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3017_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2712__S _2713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout130 input2/X vssd1 vssd1 vccd1 vccd1 _3089_/A sky130_fd_sc_hd__buf_8
XANTENNA__2849__A0 _2111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1998__S _2053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2622__S _2629_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3019__A _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ _3469_/Q _3468_/Q _3467_/Q _2250_/D vssd1 vssd1 vccd1 vccd1 _2250_/X sky130_fd_sc_hd__or4_1
XFILLER_0_18_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2181_ _3491_/Q _2587_/C _2214_/A vssd1 vssd1 vccd1 vccd1 _2181_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1965_ _1985_/S _1960_/X _1964_/X vssd1 vssd1 vccd1 vccd1 _1966_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1896_ _1902_/A _3523_/Q _2905_/B vssd1 vssd1 vccd1 vccd1 _1945_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3635_ _3637_/CLK hold42/X _3126_/Y vssd1 vssd1 vccd1 vccd1 _3635_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout106_A hold126/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3566_ _3571_/CLK _3566_/D _3060_/Y vssd1 vssd1 vccd1 vccd1 _3566_/Q sky130_fd_sc_hd__dfstp_1
X_2517_ _2516_/X _2515_/X _2551_/S vssd1 vssd1 vccd1 vccd1 _2517_/X sky130_fd_sc_hd__mux2_1
X_3497_ _3499_/CLK _3497_/D _2991_/Y vssd1 vssd1 vccd1 vccd1 _3497_/Q sky130_fd_sc_hd__dfrtp_1
X_2448_ _3402_/Q _3393_/Q _3384_/Q _3429_/Q _1943_/B _1942_/A vssd1 vssd1 vccd1 vccd1
+ _2448_/X sky130_fd_sc_hd__mux4_1
X_2379_ _2378_/X _2145_/A _2379_/S vssd1 vssd1 vccd1 vccd1 _3348_/D sky130_fd_sc_hd__mux2_1
XANTENNA__2707__S _2713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1968__S1 _2044_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2298__A1 hold14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2617__S _2618_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1750_ hold983/X _2383_/C _1749_/X vssd1 vssd1 vccd1 vccd1 _1750_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_80_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1681_ _3605_/Q hold14/X hold21/X vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__mux2_1
XFILLER_0_20_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold408 _3258_/Q vssd1 vssd1 vccd1 vccd1 hold408/X sky130_fd_sc_hd__dlygate4sd3_1
X_3420_ _3582_/CLK _3420_/D vssd1 vssd1 vccd1 vccd1 _3420_/Q sky130_fd_sc_hd__dfxtp_1
Xhold419 _2813_/X vssd1 vssd1 vccd1 vccd1 _3331_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3351_ _3369_/CLK _3351_/D vssd1 vssd1 vccd1 vccd1 _3351_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1959__S1 _2044_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2302_ hold72/X hold33/X hold30/X vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__mux2_1
XFILLER_0_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _3325_/CLK _3282_/D vssd1 vssd1 vccd1 vccd1 _3282_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2233_ _2261_/B _2238_/A vssd1 vssd1 vccd1 vccd1 _2236_/A sky130_fd_sc_hd__nand2_1
X_2164_ _3525_/Q _2164_/B vssd1 vssd1 vccd1 vccd1 _2165_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_45_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2095_ _2108_/B _2094_/X _2108_/A vssd1 vssd1 vccd1 vccd1 _2095_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2997_ _3121_/A vssd1 vssd1 vccd1 vccd1 _2997_/Y sky130_fd_sc_hd__inv_2
X_1948_ _3522_/Q _1893_/Y _1931_/B _1944_/Y _1947_/Y vssd1 vssd1 vccd1 vccd1 _1948_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_43_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1879_ _1879_/A _1879_/B vssd1 vssd1 vccd1 vccd1 _1879_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold931 _3531_/Q vssd1 vssd1 vccd1 vccd1 _1877_/A sky130_fd_sc_hd__buf_1
Xhold920 _3539_/Q vssd1 vssd1 vccd1 vccd1 _1583_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3618_ _3629_/CLK _3618_/D _3109_/Y vssd1 vssd1 vccd1 vccd1 _3618_/Q sky130_fd_sc_hd__dfrtp_1
Xhold942 _3460_/Q vssd1 vssd1 vccd1 vccd1 _2272_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 _3562_/Q vssd1 vssd1 vccd1 vccd1 _1763_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 _2157_/X vssd1 vssd1 vccd1 vccd1 _3498_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 _3528_/Q vssd1 vssd1 vccd1 vccd1 _1883_/A sky130_fd_sc_hd__buf_1
Xhold997 _1740_/X vssd1 vssd1 vccd1 vccd1 _1741_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3549_ _3559_/CLK _3549_/D _3043_/Y vssd1 vssd1 vccd1 vccd1 _3549_/Q sky130_fd_sc_hd__dfrtp_1
Xhold975 _3565_/Q vssd1 vssd1 vccd1 vccd1 hold975/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2900__S _2904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2920_ _3055_/A vssd1 vssd1 vccd1 vccd1 _2920_/Y sky130_fd_sc_hd__inv_2
X_2851_ _2074_/X hold764/X _2853_/S vssd1 vssd1 vccd1 vccd1 _2851_/X sky130_fd_sc_hd__mux2_1
X_2782_ _2812_/A1 hold278/X _2783_/S vssd1 vssd1 vccd1 vccd1 _2782_/X sky130_fd_sc_hd__mux2_1
X_1802_ _1802_/A _1802_/B vssd1 vssd1 vccd1 vccd1 _3558_/D sky130_fd_sc_hd__and2_1
XFILLER_0_86_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1733_ _3534_/Q _1596_/Y _1721_/Y _1729_/Y _1730_/Y vssd1 vssd1 vccd1 vccd1 _1735_/C
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2810__S _2813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold216 _3612_/Q vssd1 vssd1 vccd1 vccd1 _1574_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 _3640_/Q vssd1 vssd1 vccd1 vccd1 _1558_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 _2747_/X vssd1 vssd1 vccd1 vccd1 _3271_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3403_ _3403_/CLK _3403_/D vssd1 vssd1 vccd1 vccd1 _3403_/Q sky130_fd_sc_hd__dfxtp_1
Xhold227 _3235_/Q vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
X_1664_ _3614_/Q _2397_/A _1667_/S vssd1 vssd1 vccd1 vccd1 _1664_/X sky130_fd_sc_hd__mux2_1
Xhold249 _2807_/X vssd1 vssd1 vccd1 vccd1 _3325_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1595_ hold98/X vssd1 vssd1 vccd1 vccd1 _1595_/Y sky130_fd_sc_hd__inv_2
X_3334_ _3414_/CLK _3334_/D vssd1 vssd1 vccd1 vccd1 _3334_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _3305_/CLK _3265_/D vssd1 vssd1 vccd1 vccd1 _3265_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ _2216_/A _2216_/B vssd1 vssd1 vccd1 vccd1 _2216_/X sky130_fd_sc_hd__or2_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ _3403_/CLK _3196_/D vssd1 vssd1 vccd1 vccd1 _3196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2682__A1 _2813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2147_ _2156_/A _2160_/B vssd1 vssd1 vccd1 vccd1 _2147_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_72_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2078_ _2073_/X _2077_/Y _2075_/Y vssd1 vssd1 vccd1 vccd1 _2079_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_63_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold750 _3175_/Q vssd1 vssd1 vccd1 vccd1 hold750/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold761 _2612_/X vssd1 vssd1 vccd1 vccd1 _3154_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 _3185_/Q vssd1 vssd1 vccd1 vccd1 hold772/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 _3390_/Q vssd1 vssd1 vccd1 vccd1 hold794/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 _2881_/X vssd1 vssd1 vccd1 vccd1 _3406_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2036__S0 _1590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3050_ _3070_/A vssd1 vssd1 vccd1 vccd1 _3050_/Y sky130_fd_sc_hd__inv_2
X_2001_ _1999_/X _2000_/X _2045_/S vssd1 vssd1 vccd1 vccd1 _2001_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2805__S _2813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2903_ hold616/X _2076_/X _2904_/S vssd1 vssd1 vccd1 vccd1 _2903_/X sky130_fd_sc_hd__mux2_1
X_2834_ _2885_/C _3526_/Q _3525_/Q vssd1 vssd1 vccd1 vccd1 _2843_/S sky130_fd_sc_hd__or3b_4
XFILLER_0_45_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2765_ _2805_/A1 hold265/X _2773_/S vssd1 vssd1 vccd1 vccd1 _2765_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1945__A _2551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1716_ _3444_/Q _3527_/Q vssd1 vssd1 vccd1 vccd1 _1716_/X sky130_fd_sc_hd__and2b_1
X_2696_ _2806_/A1 hold152/X _2703_/S vssd1 vssd1 vccd1 vccd1 _2696_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1647_ _2393_/A hold59/X vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__nor2_1
X_1578_ _3608_/Q vssd1 vssd1 vccd1 vccd1 _1578_/Y sky130_fd_sc_hd__inv_2
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3317_ _3318_/CLK _3317_/D vssd1 vssd1 vccd1 vccd1 _3317_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _3488_/CLK _3248_/D vssd1 vssd1 vccd1 vccd1 _3248_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3179_ _3403_/CLK _3179_/D vssd1 vssd1 vccd1 vccd1 _3179_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2502__S1 _2550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2450__S _2551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold580 _3355_/Q vssd1 vssd1 vccd1 vccd1 hold580/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold591 _2624_/X vssd1 vssd1 vccd1 vccd1 _3164_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1590__A _1590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2625__S _2629_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2550_ _3187_/Q _3340_/Q _3169_/Q _3151_/Q _1911_/C _2550_/S1 vssd1 vssd1 vccd1 vccd1
+ _2550_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2582__B1 _2583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2481_ _3627_/Q hold7/A _2474_/X _2480_/X hold96/A vssd1 vssd1 vccd1 vccd1 _2481_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_50_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3102_ _3105_/A vssd1 vssd1 vccd1 vccd1 _3102_/Y sky130_fd_sc_hd__inv_2
X_3033_ _3036_/A vssd1 vssd1 vccd1 vccd1 _3033_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_85_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2817_ hold542/X _2105_/A _2823_/S vssd1 vssd1 vccd1 vccd1 _2817_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2748_ _2808_/A1 hold144/X _2753_/S vssd1 vssd1 vccd1 vccd1 _2748_/X sky130_fd_sc_hd__mux2_1
X_2679_ hold321/X _2810_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2679_/X sky130_fd_sc_hd__mux2_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2487__S0 _2554_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2800__A1 _2810_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2316__B1 _2029_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2867__A1 _2097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1981_ _1979_/X _1980_/X _2045_/S vssd1 vssd1 vccd1 vccd1 _1981_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3651_ _3659_/A vssd1 vssd1 vccd1 vccd1 _3651_/X sky130_fd_sc_hd__buf_1
X_2602_ _2105_/A hold712/X _2608_/S vssd1 vssd1 vccd1 vccd1 _2602_/X sky130_fd_sc_hd__mux2_1
X_3582_ _3582_/CLK input1/X vssd1 vssd1 vccd1 vccd1 _3582_/Q sky130_fd_sc_hd__dfxtp_1
X_2533_ _2532_/X _2531_/X _2551_/S vssd1 vssd1 vccd1 vccd1 _2533_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2464_ _3626_/Q hold7/A _2463_/X hold96/A vssd1 vssd1 vccd1 vccd1 _2464_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2395_ _2395_/A _2403_/B vssd1 vssd1 vccd1 vccd1 _3585_/D sky130_fd_sc_hd__and2_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3016_ _3114_/A vssd1 vssd1 vccd1 vccd1 _3016_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2469__S0 _2554_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout120 _3089_/A vssd1 vssd1 vccd1 vccd1 _3121_/A sky130_fd_sc_hd__buf_6
XANTENNA__3125__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2785__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2903__S _2904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2180_ _2214_/A _2180_/B _2804_/A vssd1 vssd1 vccd1 vccd1 _2180_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_75_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2776__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2813__S _2813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1964_ _1985_/S _1964_/B vssd1 vssd1 vccd1 vccd1 _1964_/X sky130_fd_sc_hd__and2b_1
XANTENNA__2240__A2 _1889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3634_ _3637_/CLK hold9/X _3125_/Y vssd1 vssd1 vccd1 vccd1 _3634_/Q sky130_fd_sc_hd__dfstp_1
X_1895_ _1933_/A _1895_/B vssd1 vssd1 vccd1 vccd1 _3526_/D sky130_fd_sc_hd__nor2_1
X_3565_ _3580_/CLK _3565_/D _3059_/Y vssd1 vssd1 vccd1 vccd1 _3565_/Q sky130_fd_sc_hd__dfstp_1
X_2516_ _3184_/Q _3337_/Q _3166_/Q _3148_/Q _1943_/B _2550_/S1 vssd1 vssd1 vccd1 vccd1
+ _2516_/X sky130_fd_sc_hd__mux4_1
X_3496_ _3499_/CLK _3496_/D _2990_/Y vssd1 vssd1 vccd1 vccd1 _3496_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2447_ _3445_/Q hold29/A _2436_/X _2446_/X _2583_/B vssd1 vssd1 vccd1 vccd1 _2447_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2700__A0 _2810_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2378_ _2383_/A _2378_/B vssd1 vssd1 vccd1 vccd1 _2378_/X sky130_fd_sc_hd__and2_1
XFILLER_0_78_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2767__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2633__S _2640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold409 _2732_/X vssd1 vssd1 vccd1 vccd1 _3258_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1680_ _2393_/A hold20/X vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__nor2_1
X_3350_ _3403_/CLK _3350_/D vssd1 vssd1 vccd1 vccd1 _3350_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2301_ _1720_/B hold52/X hold30/X vssd1 vssd1 vccd1 vccd1 _2301_/X sky130_fd_sc_hd__mux2_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _3325_/CLK _3281_/D vssd1 vssd1 vccd1 vccd1 _3281_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2232_ _2260_/A _2260_/B _2241_/A vssd1 vssd1 vccd1 vccd1 _2238_/A sky130_fd_sc_hd__and3_1
XANTENNA__2808__S _2813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2163_ _3526_/Q _2163_/B vssd1 vssd1 vccd1 vccd1 _2163_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_24_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2094_ _1581_/Y _2084_/B _2085_/Y _2089_/Y _3625_/Q _2071_/A vssd1 vssd1 vccd1 vccd1
+ _2094_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2543__S _2551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2996_ _3121_/A vssd1 vssd1 vccd1 vccd1 _2996_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2749__A0 _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1947_ _3522_/Q _1893_/Y _1945_/X _1946_/Y vssd1 vssd1 vccd1 vccd1 _1947_/Y sky130_fd_sc_hd__o211ai_1
X_1878_ _1835_/A _1840_/Y _1877_/X _1877_/A _1560_/Y vssd1 vssd1 vccd1 vccd1 _1878_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_31_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold921 _1862_/X vssd1 vssd1 vccd1 vccd1 _3539_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3617_ _3631_/CLK _3617_/D _3108_/Y vssd1 vssd1 vccd1 vccd1 _3617_/Q sky130_fd_sc_hd__dfrtp_1
Xhold910 _2355_/X vssd1 vssd1 vccd1 vccd1 _3343_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 _1878_/X vssd1 vssd1 vccd1 vccd1 _3531_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 _2286_/X vssd1 vssd1 vccd1 vccd1 _3460_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3548_ _3576_/CLK _3548_/D _3042_/Y vssd1 vssd1 vccd1 vccd1 _3548_/Q sky130_fd_sc_hd__dfrtp_1
Xhold954 _3526_/Q vssd1 vssd1 vccd1 vccd1 _1893_/A sky130_fd_sc_hd__buf_1
Xhold987 _1884_/X vssd1 vssd1 vccd1 vccd1 _3528_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 _1741_/Y vssd1 vssd1 vccd1 vccd1 wire80/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 _1766_/X vssd1 vssd1 vccd1 vccd1 _3562_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 _1760_/X vssd1 vssd1 vccd1 vccd1 _3565_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3479_ _3499_/CLK _3479_/D _2973_/Y vssd1 vssd1 vccd1 vccd1 _3479_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2453__S _2551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2912__A0 _2075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2628__S _2629_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2850_ _2067_/Y hold752/X _2853_/S vssd1 vssd1 vccd1 vccd1 _2850_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1801_ _1797_/B _1803_/A _1803_/B _1797_/A vssd1 vssd1 vccd1 vccd1 _1802_/B sky130_fd_sc_hd__a31o_1
X_2781_ _2811_/A1 hold317/X _2783_/S vssd1 vssd1 vccd1 vccd1 _2781_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1732_ _3447_/Q _1879_/A _1845_/A _1595_/Y vssd1 vssd1 vccd1 vccd1 _1735_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_25_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold217 _3244_/Q vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
X_1663_ _2585_/B _2410_/A _2419_/A vssd1 vssd1 vccd1 vccd1 _1663_/X sky130_fd_sc_hd__and3_1
Xhold206 _3639_/Q vssd1 vssd1 vccd1 vccd1 _1559_/A sky130_fd_sc_hd__dlygate4sd3_1
X_3402_ _3414_/CLK _3402_/D vssd1 vssd1 vccd1 vccd1 _3402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold228 _2707_/X vssd1 vssd1 vccd1 vccd1 _3235_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 _3197_/Q vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
X_1594_ _3458_/Q vssd1 vssd1 vccd1 vccd1 _2580_/A sky130_fd_sc_hd__inv_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _3414_/CLK _3333_/D vssd1 vssd1 vccd1 vccd1 _3333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2111__B _2111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _3318_/CLK _3264_/D vssd1 vssd1 vccd1 vccd1 _3264_/Q sky130_fd_sc_hd__dfxtp_1
X_2215_ _2212_/Y _2213_/X _2214_/Y _2214_/B _2211_/A vssd1 vssd1 vccd1 vccd1 _2215_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _3369_/CLK _3195_/D vssd1 vssd1 vccd1 vccd1 _3195_/Q sky130_fd_sc_hd__dfxtp_1
X_2146_ _2149_/A _2367_/C _2149_/B vssd1 vssd1 vccd1 vccd1 _2160_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2077_ _2338_/B vssd1 vssd1 vccd1 vccd1 _2077_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_88_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2979_ _3126_/A vssd1 vssd1 vccd1 vccd1 _2979_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2198__A1 _2222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold751 _2637_/X vssd1 vssd1 vccd1 vccd1 _3175_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold740 _3417_/Q vssd1 vssd1 vccd1 vccd1 hold740/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 _3176_/Q vssd1 vssd1 vccd1 vccd1 hold762/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 _2648_/X vssd1 vssd1 vccd1 vccd1 _3185_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 _2863_/X vssd1 vssd1 vccd1 vccd1 _3390_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 _3408_/Q vssd1 vssd1 vccd1 vccd1 hold784/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_18_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3614_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2911__S _2914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2036__S1 _2222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2000_ hold362/X hold428/X hold358/X hold398/X _2044_/S0 _2044_/S1 vssd1 vssd1 vccd1
+ vccd1 _2000_/X sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2902_ hold656/X _2074_/X _2904_/S vssd1 vssd1 vccd1 vccd1 _2902_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2833_ hold520/X _2339_/B _2833_/S vssd1 vssd1 vccd1 vccd1 _2833_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2764_ _2764_/A _2794_/A _2794_/B vssd1 vssd1 vccd1 vccd1 _2773_/S sky130_fd_sc_hd__or3b_4
X_1715_ _3527_/Q _3444_/Q vssd1 vssd1 vccd1 vccd1 _1715_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2695_ _2805_/A1 hold282/X _2703_/S vssd1 vssd1 vccd1 vccd1 _2695_/X sky130_fd_sc_hd__mux2_1
X_1646_ hold58/X _1646_/B vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__or2_2
X_1577_ _3609_/Q vssd1 vssd1 vccd1 vccd1 _1577_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_6_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3316_ _3316_/CLK _3316_/D vssd1 vssd1 vccd1 vccd1 _3316_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ _3316_/CLK _3247_/D vssd1 vssd1 vccd1 vccd1 _3247_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3178_ _3427_/CLK _3178_/D vssd1 vssd1 vccd1 vccd1 _3178_/Q sky130_fd_sc_hd__dfxtp_1
X_2129_ _2129_/A _2160_/A vssd1 vssd1 vccd1 vccd1 _2130_/C sky130_fd_sc_hd__or2_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1918__A1 _1911_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2591__A1 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold581 _2830_/X vssd1 vssd1 vccd1 vccd1 _3355_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold570 _3420_/Q vssd1 vssd1 vccd1 vccd1 hold570/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 _3424_/Q vssd1 vssd1 vccd1 vccd1 hold592/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2906__S _2914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2480_ _3518_/Q _2507_/B _2475_/X _2479_/X hold59/A vssd1 vssd1 vccd1 vccd1 _2480_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_50_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3101_ _3105_/A vssd1 vssd1 vccd1 vccd1 _3101_/Y sky130_fd_sc_hd__inv_2
X_3032_ _3036_/A vssd1 vssd1 vccd1 vccd1 _3032_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_73_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1659__C input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2816_ hold552/X _2097_/A _2823_/S vssd1 vssd1 vccd1 vccd1 _2816_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2551__S _2551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout129_A _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2747_ _2807_/A1 hold237/X _2753_/S vssd1 vssd1 vccd1 vccd1 _2747_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2678_ hold428/X _2809_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2678_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1629_ hold6/X _1646_/B vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__or2_4
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2487__S1 _1911_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_33_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3563_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2636__S _2640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1980_ _3221_/Q _3212_/Q _3203_/Q _3329_/Q _2224_/B _2193_/A1 vssd1 vssd1 vccd1 vccd1
+ _1980_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_82_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3650_ _3659_/A vssd1 vssd1 vccd1 vccd1 _3650_/X sky130_fd_sc_hd__buf_1
X_2601_ _2097_/A hold788/X _2608_/S vssd1 vssd1 vccd1 vccd1 _2601_/X sky130_fd_sc_hd__mux2_1
X_3581_ _3631_/CLK _3581_/D _3074_/Y vssd1 vssd1 vccd1 vccd1 _3581_/Q sky130_fd_sc_hd__dfrtp_4
X_2532_ _3176_/Q _3425_/Q _3416_/Q _3158_/Q _2554_/S0 _1942_/A vssd1 vssd1 vccd1 vccd1
+ _2532_/X sky130_fd_sc_hd__mux4_1
XANTENNA__1989__S0 _2044_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2307__A1 _2585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2463_ _3617_/Q _1645_/Y _2461_/X _2462_/X _2571_/B vssd1 vssd1 vccd1 vccd1 _2463_/X
+ sky130_fd_sc_hd__a221o_1
X_2394_ _2585_/A _2403_/B vssd1 vssd1 vccd1 vccd1 _3584_/D sky130_fd_sc_hd__and2_1
XANTENNA__2400__A hold52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2546__S _2551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3015_ _3089_/A vssd1 vssd1 vccd1 vccd1 _3015_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2491__B1 _2483_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2469__S1 _1911_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout121 _3089_/A vssd1 vssd1 vccd1 vccd1 _3105_/A sky130_fd_sc_hd__buf_8
XFILLER_0_10_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout110 hold120/X vssd1 vssd1 vccd1 vccd1 _2806_/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_10_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2980__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output42_A _2570_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2473__B1 _2465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1963_ _1962_/X _1961_/X _2045_/S vssd1 vssd1 vccd1 vccd1 _1964_/B sky130_fd_sc_hd__mux2_1
X_1894_ _2824_/B hold955/X _2598_/C vssd1 vssd1 vccd1 vccd1 _1894_/X sky130_fd_sc_hd__mux2_1
X_3633_ _3633_/CLK hold24/X _3124_/Y vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfstp_1
XFILLER_0_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3564_ _3580_/CLK _3564_/D _3058_/Y vssd1 vssd1 vccd1 vccd1 _3564_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2515_ _3406_/Q _3397_/Q _3388_/Q _3433_/Q _1943_/B _2550_/S1 vssd1 vssd1 vccd1 vccd1
+ _2515_/X sky130_fd_sc_hd__mux4_1
X_3495_ _3623_/CLK _3495_/D _2989_/Y vssd1 vssd1 vccd1 vccd1 _3495_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2446_ _3625_/Q hold7/A _2437_/X _2445_/X hold96/A vssd1 vssd1 vccd1 vccd1 _2446_/X
+ sky130_fd_sc_hd__o221a_1
X_2377_ _3346_/Q _2366_/X _2370_/A _2145_/D _2379_/S vssd1 vssd1 vccd1 vccd1 _2377_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_78_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2455__B1 _2447_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2914__S _2914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2550__S0 _1911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2758__A1 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3280_ _3305_/CLK _3280_/D vssd1 vssd1 vccd1 vccd1 _3280_/Q sky130_fd_sc_hd__dfxtp_1
X_2300_ hold62/X hold44/X hold30/X vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__mux2_1
XFILLER_0_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ _2231_/A _2231_/B wire80/X _2231_/D vssd1 vssd1 vccd1 vccd1 _2241_/A sky130_fd_sc_hd__and4_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2162_ _3526_/Q _2163_/B vssd1 vssd1 vccd1 vccd1 _2162_/X sky130_fd_sc_hd__or2_1
X_2093_ _2060_/Y _2069_/B _2088_/B _2062_/B _2071_/A _1783_/A vssd1 vssd1 vccd1 vccd1
+ _2108_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2541__S0 _1943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2995_ _3055_/A vssd1 vssd1 vccd1 vccd1 _2995_/Y sky130_fd_sc_hd__inv_2
X_1946_ _1945_/B _1945_/C _2551_/S vssd1 vssd1 vccd1 vccd1 _1946_/Y sky130_fd_sc_hd__o21ai_1
X_1877_ _1877_/A _1877_/B vssd1 vssd1 vccd1 vccd1 _1877_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold900 _3538_/Q vssd1 vssd1 vccd1 vccd1 _1849_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 _3542_/Q vssd1 vssd1 vccd1 vccd1 _1855_/A sky130_fd_sc_hd__buf_1
Xhold922 _3467_/Q vssd1 vssd1 vccd1 vccd1 hold922/X sky130_fd_sc_hd__dlygate4sd3_1
X_3616_ _3629_/CLK _3616_/D _3107_/Y vssd1 vssd1 vccd1 vccd1 _3616_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout111_A hold120/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold933 _3534_/Q vssd1 vssd1 vccd1 vccd1 _1871_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3547_ _3576_/CLK _3547_/D _3041_/Y vssd1 vssd1 vccd1 vccd1 _3547_/Q sky130_fd_sc_hd__dfrtp_1
Xhold955 _1893_/Y vssd1 vssd1 vccd1 vccd1 hold955/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 _3568_/Q vssd1 vssd1 vccd1 vccd1 _1751_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 _3564_/Q vssd1 vssd1 vccd1 vccd1 hold977/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 _3476_/Q vssd1 vssd1 vccd1 vccd1 _1956_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold988 _3499_/Q vssd1 vssd1 vccd1 vccd1 _1589_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold999 _1950_/B vssd1 vssd1 vccd1 vccd1 _2367_/B sky130_fd_sc_hd__dlygate4sd3_1
X_3478_ _3499_/CLK _3478_/D _2972_/Y vssd1 vssd1 vccd1 vccd1 _3478_/Q sky130_fd_sc_hd__dfrtp_1
X_2429_ _3179_/Q _3332_/Q _3161_/Q _3143_/Q _1943_/B _1942_/A vssd1 vssd1 vccd1 vccd1
+ _2429_/X sky130_fd_sc_hd__mux4_1
XANTENNA__2685__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2532__S0 _2554_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2909__S _2914_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1651__A1 hold33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1800_ _1778_/A _1802_/A _1799_/X vssd1 vssd1 vccd1 vccd1 _1800_/X sky130_fd_sc_hd__a21o_1
X_2780_ _2810_/A1 hold319/X _2783_/S vssd1 vssd1 vccd1 vccd1 _2780_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1731_ _3528_/Q _3445_/Q vssd1 vssd1 vccd1 vccd1 _1731_/X sky130_fd_sc_hd__and2b_1
XANTENNA__2600__A0 _2342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1662_ _2410_/A _2407_/A vssd1 vssd1 vccd1 vccd1 _2439_/A sky130_fd_sc_hd__and2_1
Xhold207 hold207/A vssd1 vssd1 vccd1 vccd1 _1834_/A sky130_fd_sc_hd__clkbuf_2
Xhold218 _2717_/X vssd1 vssd1 vccd1 vccd1 _3244_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3401_ _3526_/CLK _3401_/D vssd1 vssd1 vccd1 vccd1 _3401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold229 _3217_/Q vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__dlygate4sd3_1
X_1593_ _3462_/Q vssd1 vssd1 vccd1 vccd1 _1593_/Y sky130_fd_sc_hd__inv_2
X_3332_ _3403_/CLK _3332_/D vssd1 vssd1 vccd1 vccd1 _3332_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _3318_/CLK _3263_/D vssd1 vssd1 vccd1 vccd1 _3263_/Q sky130_fd_sc_hd__dfxtp_1
X_2214_ _2214_/A _2214_/B vssd1 vssd1 vccd1 vccd1 _2214_/Y sky130_fd_sc_hd__nor2_1
X_3194_ _3416_/CLK _3194_/D vssd1 vssd1 vccd1 vccd1 _3194_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2667__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2145_ _2145_/A _2378_/B _3346_/Q _2145_/D vssd1 vssd1 vccd1 vccd1 _2149_/B sky130_fd_sc_hd__or4_2
XFILLER_0_88_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2076_ _2108_/A _2076_/B _2076_/C vssd1 vssd1 vccd1 vccd1 _2076_/X sky130_fd_sc_hd__and3_1
XANTENNA__1642__A1 _2396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2978_ _3126_/A vssd1 vssd1 vccd1 vccd1 _2978_/Y sky130_fd_sc_hd__inv_2
X_1929_ _1929_/A _1929_/B vssd1 vssd1 vccd1 vccd1 _1930_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_71_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold730 _3196_/Q vssd1 vssd1 vccd1 vccd1 hold730/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold752 _3373_/Q vssd1 vssd1 vccd1 vccd1 hold752/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 _2893_/X vssd1 vssd1 vccd1 vccd1 _3417_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 _2638_/X vssd1 vssd1 vccd1 vccd1 _3176_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 _3168_/Q vssd1 vssd1 vccd1 vccd1 hold796/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 _2883_/X vssd1 vssd1 vccd1 vccd1 _3408_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 _3161_/Q vssd1 vssd1 vccd1 vccd1 hold774/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1633__S hold8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2658__A0 _2075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1633__A1 hold41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2639__S _2640_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2649__A0 _2338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
X_2901_ hold592/X _2067_/Y _2904_/S vssd1 vssd1 vccd1 vccd1 _2901_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2832_ hold528/X _2338_/B _2833_/S vssd1 vssd1 vccd1 vccd1 _2832_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2763_ hold366/X _2813_/A1 _2763_/S vssd1 vssd1 vccd1 vccd1 _2763_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2403__A hold14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1714_ _3538_/Q hold46/X vssd1 vssd1 vccd1 vccd1 _1714_/Y sky130_fd_sc_hd__nand2b_1
X_2694_ _2794_/B _2804_/A _2794_/A vssd1 vssd1 vccd1 vccd1 _2703_/S sky130_fd_sc_hd__or3b_4
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1645_ hold58/A _1646_/B vssd1 vssd1 vccd1 vccd1 _1645_/Y sky130_fd_sc_hd__nor2_2
X_1576_ _3610_/Q vssd1 vssd1 vccd1 vccd1 _2476_/A sky130_fd_sc_hd__inv_2
X_3315_ _3319_/CLK _3315_/D vssd1 vssd1 vccd1 vccd1 _3315_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ _3318_/CLK _3246_/D vssd1 vssd1 vccd1 vccd1 _3246_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3177_ _3583_/CLK _3177_/D vssd1 vssd1 vccd1 vccd1 _3177_/Q sky130_fd_sc_hd__dfxtp_1
X_2128_ _2366_/B _2366_/C vssd1 vssd1 vccd1 vccd1 _2133_/B sky130_fd_sc_hd__nand2_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2059_ _2059_/A _2089_/B vssd1 vssd1 vccd1 vccd1 _2067_/B sky130_fd_sc_hd__nand2_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1918__A2 _2554_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2879__A0 _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold571 _2897_/X vssd1 vssd1 vccd1 vccd1 _3420_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold560 _3407_/Q vssd1 vssd1 vccd1 vccd1 hold560/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 _2901_/X vssd1 vssd1 vccd1 vccd1 _3424_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 _3401_/Q vssd1 vssd1 vccd1 vccd1 hold582/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2343__A2 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2983__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1599__A _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2334__A2 _1889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3100_ _3126_/A vssd1 vssd1 vccd1 vccd1 _3100_/Y sky130_fd_sc_hd__inv_2
X_3031_ _3128_/A vssd1 vssd1 vccd1 vccd1 _3031_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_3_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3331_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2270__A1 _1889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2815_ hold554/X _2342_/B _2823_/S vssd1 vssd1 vccd1 vccd1 _2815_/X sky130_fd_sc_hd__mux2_1
X_2746_ _2806_/A1 hold173/X _2753_/S vssd1 vssd1 vccd1 vccd1 _2746_/X sky130_fd_sc_hd__mux2_1
X_2677_ hold142/X _2808_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2677_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1628_ hold6/A _1646_/B vssd1 vssd1 vccd1 vccd1 _2571_/B sky130_fd_sc_hd__nor2_2
X_1559_ _1559_/A vssd1 vssd1 vccd1 vccd1 _2367_/A sky130_fd_sc_hd__inv_2
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3229_ _3325_/CLK _3229_/D vssd1 vssd1 vccd1 vccd1 _3229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1964__A_N _1985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2978__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold390 _3284_/Q vssd1 vssd1 vccd1 vccd1 hold390/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2600_ _2342_/B hold710/X _2608_/S vssd1 vssd1 vccd1 vccd1 _2600_/X sky130_fd_sc_hd__mux2_1
X_3580_ _3580_/CLK _3580_/D vssd1 vssd1 vccd1 vccd1 _3580_/Q sky130_fd_sc_hd__dfxtp_1
X_2531_ _3374_/Q _3356_/Q _3365_/Q _3194_/Q _2554_/S0 _1942_/A vssd1 vssd1 vccd1 vccd1
+ _2531_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_23_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1989__S1 _2044_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2462_ _3517_/Q _2507_/B hold59/A vssd1 vssd1 vccd1 vccd1 _2462_/X sky130_fd_sc_hd__o21a_1
X_2393_ _2393_/A hold67/X vssd1 vssd1 vccd1 vccd1 _2403_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_3_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3014_ _3089_/A vssd1 vssd1 vccd1 vccd1 _3014_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2491__A1 _2506_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2729_ _2809_/A1 hold392/X _2733_/S vssd1 vssd1 vccd1 vccd1 _2729_/X sky130_fd_sc_hd__mux2_1
Xfanout100 hold927/X vssd1 vssd1 vccd1 vccd1 _1811_/A sky130_fd_sc_hd__buf_4
Xfanout111 hold120/X vssd1 vssd1 vccd1 vccd1 _2395_/A sky130_fd_sc_hd__clkbuf_4
Xfanout122 _3089_/A vssd1 vssd1 vccd1 vccd1 _3095_/A sky130_fd_sc_hd__buf_4
XANTENNA__1641__S hold8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2472__S _3522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2473__A1 _2506_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1962_ hold459/X hold463/X hold349/X hold378/X _1590_/A _2193_/A1 vssd1 vssd1 vccd1
+ vccd1 _1962_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_83_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1893_ _1893_/A _1945_/B vssd1 vssd1 vccd1 vccd1 _1893_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3632_ _3637_/CLK hold55/X _3123_/Y vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__dfstp_1
XFILLER_0_70_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3563_ _3563_/CLK _3563_/D _3057_/Y vssd1 vssd1 vccd1 vccd1 _3563_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2514_ _2510_/X _2511_/Y _2513_/X _2511_/B hold72/A vssd1 vssd1 vccd1 vccd1 _2514_/X
+ sky130_fd_sc_hd__a32o_1
X_3494_ _3610_/CLK _3494_/D _2988_/Y vssd1 vssd1 vccd1 vccd1 _3494_/Q sky130_fd_sc_hd__dfrtp_1
X_2445_ _3516_/Q _2507_/B _2438_/X _2444_/X hold59/A vssd1 vssd1 vccd1 vccd1 _2445_/X
+ sky130_fd_sc_hd__o221a_1
X_2376_ _1824_/A _1793_/A _2370_/A _1808_/D _1772_/B vssd1 vssd1 vccd1 vccd1 _2376_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_78_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1636__S hold8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2040__B _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2455__A1 _2506_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2991__A _3131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2550__S1 _2550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2038__A_N _1985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ hold476/X _2229_/X _2188_/Y vssd1 vssd1 vccd1 vccd1 _2230_/X sky130_fd_sc_hd__o21a_1
X_2161_ _2160_/Y _2160_/A _2161_/S vssd1 vssd1 vccd1 vccd1 _2161_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2092_ _2097_/A vssd1 vssd1 vccd1 vccd1 _2092_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2541__S1 _2550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2994_ _3055_/A vssd1 vssd1 vccd1 vccd1 _2994_/Y sky130_fd_sc_hd__inv_2
X_1945_ _2551_/S _1945_/B _1945_/C vssd1 vssd1 vccd1 vccd1 _1945_/X sky130_fd_sc_hd__or3_1
XFILLER_0_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1876_ _1835_/A _1842_/Y _1875_/X _1841_/A _1560_/Y vssd1 vssd1 vccd1 vccd1 _1876_/X
+ sky130_fd_sc_hd__a32o_1
Xhold901 _1864_/X vssd1 vssd1 vccd1 vccd1 _3538_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 _1856_/X vssd1 vssd1 vccd1 vccd1 _3542_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3615_ _3623_/CLK _3615_/D _3106_/Y vssd1 vssd1 vccd1 vccd1 _3615_/Q sky130_fd_sc_hd__dfrtp_1
Xhold934 _1872_/X vssd1 vssd1 vccd1 vccd1 _3534_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 _3537_/Q vssd1 vssd1 vccd1 vccd1 _1865_/A sky130_fd_sc_hd__buf_1
X_3546_ _3576_/CLK _3546_/D _3040_/Y vssd1 vssd1 vccd1 vccd1 _3546_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout104_A hold33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold945 _1754_/X vssd1 vssd1 vccd1 vccd1 _3568_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 _1894_/X vssd1 vssd1 vccd1 vccd1 _1895_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 _1762_/X vssd1 vssd1 vccd1 vccd1 _3564_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 _3567_/Q vssd1 vssd1 vccd1 vccd1 hold967/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2382__B1 _1889_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold989 _2153_/X vssd1 vssd1 vccd1 vccd1 hold989/X sky130_fd_sc_hd__dlygate4sd3_1
X_3477_ _3499_/CLK _3477_/D _2971_/Y vssd1 vssd1 vccd1 vccd1 _3477_/Q sky130_fd_sc_hd__dfrtp_1
X_2428_ _3401_/Q _3392_/Q _3383_/Q _3428_/Q _1943_/B _1942_/A vssd1 vssd1 vccd1 vccd1
+ _2428_/X sky130_fd_sc_hd__mux4_1
X_2359_ _2476_/A _2211_/A _2357_/X _2358_/X hold476/X vssd1 vssd1 vccd1 vccd1 _2359_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2532__S1 _1942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2750__S _2753_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2676__A1 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1730_ _3454_/Q _1865_/A vssd1 vssd1 vccd1 vccd1 _1730_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_25_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1661_ hold65/X _1661_/B _1661_/C vssd1 vssd1 vccd1 vccd1 _2407_/A sky130_fd_sc_hd__and3b_1
Xhold208 hold208/A vssd1 vssd1 vccd1 vccd1 _1770_/S sky130_fd_sc_hd__buf_1
Xhold219 _3289_/Q vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__dlygate4sd3_1
X_3400_ _3436_/CLK _3400_/D vssd1 vssd1 vccd1 vccd1 _3400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1592_ _1592_/A vssd1 vssd1 vccd1 vccd1 _2275_/A sky130_fd_sc_hd__inv_2
XFILLER_0_21_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3331_ _3331_/CLK _3331_/D vssd1 vssd1 vccd1 vccd1 _3331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3305_/CLK _3262_/D vssd1 vssd1 vccd1 vccd1 _3262_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ _2212_/C _2212_/B _2211_/X vssd1 vssd1 vccd1 vccd1 _2213_/X sky130_fd_sc_hd__a21bo_1
X_3193_ _3416_/CLK _3193_/D vssd1 vssd1 vccd1 vccd1 _3193_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2144_ _2134_/C _2136_/C _2143_/Y vssd1 vssd1 vccd1 vccd1 _2144_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2075_ _2076_/C _2075_/B vssd1 vssd1 vccd1 vccd1 _2075_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_48_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2977_ _3126_/A vssd1 vssd1 vccd1 vccd1 _2977_/Y sky130_fd_sc_hd__inv_2
X_1928_ _1928_/A _1931_/B vssd1 vssd1 vccd1 vccd1 _1929_/B sky130_fd_sc_hd__nor2_1
X_1859_ _1859_/A _1859_/B vssd1 vssd1 vccd1 vccd1 _1859_/X sky130_fd_sc_hd__or2_1
Xhold720 _3165_/Q vssd1 vssd1 vccd1 vccd1 hold720/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 _2850_/X vssd1 vssd1 vccd1 vccd1 _3373_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 _3429_/Q vssd1 vssd1 vccd1 vccd1 hold742/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 _3374_/Q vssd1 vssd1 vccd1 vccd1 hold764/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 _2660_/X vssd1 vssd1 vccd1 vccd1 _3196_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3529_ _3542_/CLK _3529_/D _3023_/Y vssd1 vssd1 vccd1 vccd1 _3529_/Q sky130_fd_sc_hd__dfrtp_1
Xhold786 _3157_/Q vssd1 vssd1 vccd1 vccd1 hold786/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 _2628_/X vssd1 vssd1 vccd1 vccd1 _3168_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 _2621_/X vssd1 vssd1 vccd1 vccd1 _3161_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2745__S _2753_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2830__A1 _2079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3571_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2346__B1 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__clkbuf_2
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2900_ hold564/X _2109_/X _2904_/S vssd1 vssd1 vccd1 vccd1 _2900_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2821__A1 _2075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2831_ hold562/X _2075_/B _2833_/S vssd1 vssd1 vccd1 vccd1 _2831_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2762_ hold300/X _2812_/A1 _2763_/S vssd1 vssd1 vccd1 vccd1 _2762_/X sky130_fd_sc_hd__mux2_1
X_1713_ _3450_/Q _1843_/A vssd1 vssd1 vccd1 vccd1 _1713_/Y sky130_fd_sc_hd__nand2b_1
X_2693_ _2813_/A1 hold457/X _2693_/S vssd1 vssd1 vccd1 vccd1 _2693_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1644_ _2121_/A _2585_/A hold8/X vssd1 vssd1 vccd1 vccd1 _1644_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2432__S0 _1911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1575_ _1575_/A vssd1 vssd1 vccd1 vccd1 _1575_/Y sky130_fd_sc_hd__inv_2
X_3314_ _3316_/CLK _3314_/D vssd1 vssd1 vccd1 vccd1 _3314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _3318_/CLK _3245_/D vssd1 vssd1 vccd1 vccd1 _3245_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3176_ _3583_/CLK _3176_/D vssd1 vssd1 vccd1 vccd1 _3176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2127_ _2127_/A _2127_/B _2127_/C _2127_/D vssd1 vssd1 vccd1 vccd1 _2366_/C sky130_fd_sc_hd__and4_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2058_ _2059_/A _2089_/B vssd1 vssd1 vccd1 vccd1 _2076_/B sky130_fd_sc_hd__and2_1
XFILLER_0_88_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2499__S0 _1943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2812__A1 _2812_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold550 _3335_/Q vssd1 vssd1 vccd1 vccd1 hold550/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 _3190_/Q vssd1 vssd1 vccd1 vccd1 hold572/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 _2882_/X vssd1 vssd1 vccd1 vccd1 _3407_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1644__S hold8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold594 _3399_/Q vssd1 vssd1 vccd1 vccd1 hold594/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 _2876_/X vssd1 vssd1 vccd1 vccd1 _3401_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout84_A _1942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2803__A1 _2813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2223__B _2224_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3030_ _3128_/A vssd1 vssd1 vccd1 vccd1 _3030_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_53_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2814_ _2824_/B _2905_/B _2895_/C vssd1 vssd1 vccd1 vccd1 _2823_/S sky130_fd_sc_hd__nor3_4
XFILLER_0_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2745_ _2805_/A1 hold263/X _2753_/S vssd1 vssd1 vccd1 vccd1 _2745_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2676_ hold257/X _2807_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2676_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1627_ hold28/X _1668_/A vssd1 vssd1 vccd1 vccd1 _1646_/B sky130_fd_sc_hd__nand2_2
XANTENNA__2730__A0 _2810_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1558_ _1558_/A vssd1 vssd1 vccd1 vccd1 _1743_/A sky130_fd_sc_hd__inv_2
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3228_ _3331_/CLK _3228_/D vssd1 vssd1 vccd1 vccd1 _3228_/Q sky130_fd_sc_hd__dfxtp_1
X_3159_ _3583_/CLK _3159_/D vssd1 vssd1 vccd1 vccd1 _3159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1639__S hold8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold380 _3277_/Q vssd1 vssd1 vccd1 vccd1 hold380/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2721__A0 _2811_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold391 _2761_/X vssd1 vssd1 vccd1 vccd1 _3284_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_42_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3623_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2788__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2530_ _2529_/X _2528_/X _2551_/S vssd1 vssd1 vccd1 vccd1 _2530_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2461_ _3613_/Q _2439_/A _2459_/X _2460_/X _2406_/X vssd1 vssd1 vccd1 vccd1 _2461_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2712__A0 _2812_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2392_ hold95/A hold66/X vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__nand2_4
XFILLER_0_3_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3013_ _3114_/A vssd1 vssd1 vccd1 vccd1 _3013_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2779__A0 _2809_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2728_ _2808_/A1 hold128/X _2733_/S vssd1 vssd1 vccd1 vccd1 _2728_/X sky130_fd_sc_hd__mux2_1
X_2659_ _2338_/B hold644/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2659_/X sky130_fd_sc_hd__mux2_1
Xfanout112 hold176/X vssd1 vssd1 vccd1 vccd1 _2805_/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout101 hold49/X vssd1 vssd1 vccd1 vccd1 _2813_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__2703__A0 _2813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout123 _3126_/A vssd1 vssd1 vccd1 vccd1 _3124_/A sky130_fd_sc_hd__buf_8
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2753__S _2753_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1961_ hold461/X _3286_/Q _3277_/Q _3268_/Q _1590_/A _2193_/A1 vssd1 vssd1 vccd1
+ vccd1 _1961_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_28_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1892_ _2905_/B _1902_/A _3523_/Q vssd1 vssd1 vccd1 vccd1 _1945_/B sky130_fd_sc_hd__and3_1
X_3631_ _3631_/CLK hold71/X _3122_/Y vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3562_ _3563_/CLK _3562_/D _3056_/Y vssd1 vssd1 vccd1 vccd1 _3562_/Q sky130_fd_sc_hd__dfstp_1
X_2513_ _3620_/Q _1645_/Y _2568_/D _2512_/X vssd1 vssd1 vccd1 vccd1 _2513_/X sky130_fd_sc_hd__a22o_1
X_3493_ _3493_/CLK _3493_/D _2987_/Y vssd1 vssd1 vccd1 vccd1 _3493_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2444_ _3484_/Q _2507_/C _2508_/A _2443_/X vssd1 vssd1 vccd1 vccd1 _2444_/X sky130_fd_sc_hd__o211a_1
X_2375_ _2375_/A _2375_/B vssd1 vssd1 vccd1 vccd1 _3344_/D sky130_fd_sc_hd__nand2_1
XANTENNA__1672__A0 _2397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1975__A1 _1985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2748__S _2753_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ _2160_/A _2160_/B vssd1 vssd1 vccd1 vccd1 _2160_/Y sky130_fd_sc_hd__nor2_1
X_2091_ _2056_/B _2090_/X _2086_/X _2082_/Y _2076_/B vssd1 vssd1 vccd1 vccd1 _2091_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_88_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2993_ _3131_/A vssd1 vssd1 vccd1 vccd1 _2993_/Y sky130_fd_sc_hd__inv_2
X_1944_ _2165_/B _1944_/B vssd1 vssd1 vccd1 vccd1 _1944_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_83_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1957__A1 _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1875_ _1877_/A _1877_/B _1841_/A vssd1 vssd1 vccd1 vccd1 _1875_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_43_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3614_ _3614_/CLK _3614_/D _3105_/Y vssd1 vssd1 vccd1 vccd1 _3614_/Q sky130_fd_sc_hd__dfrtp_1
Xhold902 _3575_/Q vssd1 vssd1 vccd1 vccd1 _1705_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 _3573_/Q vssd1 vssd1 vccd1 vccd1 _1692_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2906__A0 _2342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold924 _1866_/X vssd1 vssd1 vccd1 vccd1 _3537_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 _3532_/Q vssd1 vssd1 vccd1 vccd1 _1841_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3545_ _3583_/CLK _3545_/D _3039_/Y vssd1 vssd1 vccd1 vccd1 _3545_/Q sky130_fd_sc_hd__dfrtp_1
Xhold946 _3524_/Q vssd1 vssd1 vccd1 vccd1 _1902_/A sky130_fd_sc_hd__buf_1
Xhold979 _3556_/Q vssd1 vssd1 vccd1 vccd1 _1803_/A sky130_fd_sc_hd__buf_1
Xhold957 _3560_/Q vssd1 vssd1 vccd1 vccd1 _1767_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 _1756_/X vssd1 vssd1 vccd1 vccd1 _3567_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3476_ _3610_/CLK _3476_/D _2970_/Y vssd1 vssd1 vccd1 vccd1 _3476_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_86_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2427_ _3444_/Q hold29/A _2583_/B _2426_/X vssd1 vssd1 vccd1 vccd1 _2427_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_86_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2358_ _2476_/A _2211_/A _2208_/A _1577_/Y vssd1 vssd1 vccd1 vccd1 _2358_/X sky130_fd_sc_hd__o22a_1
X_2289_ hold28/A _2419_/B vssd1 vssd1 vccd1 vccd1 _2511_/B sky130_fd_sc_hd__and2_4
XANTENNA__1948__A1 _3522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1890__B _2231_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2005__A_N _1985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1660_ _1660_/A input4/X input5/X input6/X vssd1 vssd1 vccd1 vccd1 _1661_/C sky130_fd_sc_hd__and4_1
Xhold209 _3618_/Q vssd1 vssd1 vccd1 vccd1 _1570_/A sky130_fd_sc_hd__dlygate4sd3_1
X_1591_ _1956_/A vssd1 vssd1 vccd1 vccd1 _2187_/A sky130_fd_sc_hd__inv_2
XFILLER_0_0_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3330_ _3330_/CLK _3330_/D vssd1 vssd1 vccd1 vccd1 _3330_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _3319_/CLK _3261_/D vssd1 vssd1 vccd1 vccd1 _3261_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ _2211_/X _2212_/B _2212_/C vssd1 vssd1 vccd1 vccd1 _2212_/Y sky130_fd_sc_hd__nand3b_1
X_3192_ _3414_/CLK _3192_/D vssd1 vssd1 vccd1 vccd1 _3192_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2143_ _2130_/A _2136_/C _2134_/C vssd1 vssd1 vccd1 vccd1 _2143_/Y sky130_fd_sc_hd__a21oi_1
X_2074_ _2080_/A _2070_/X _2072_/Y _2108_/A _2076_/B vssd1 vssd1 vccd1 vccd1 _2074_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_88_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2136__B _3346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2976_ _3105_/A vssd1 vssd1 vccd1 vccd1 _2976_/Y sky130_fd_sc_hd__inv_2
X_1927_ _2350_/B _1931_/B _1926_/Y vssd1 vssd1 vccd1 vccd1 _1930_/A sky130_fd_sc_hd__a21bo_1
X_1858_ _1858_/A _1858_/B vssd1 vssd1 vccd1 vccd1 _3541_/D sky130_fd_sc_hd__and2_1
XFILLER_0_16_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold721 _2625_/X vssd1 vssd1 vccd1 vccd1 _3165_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold710 _3143_/Q vssd1 vssd1 vccd1 vccd1 hold710/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold743 _2907_/X vssd1 vssd1 vccd1 vccd1 _3429_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 _3148_/Q vssd1 vssd1 vccd1 vccd1 hold754/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 _3194_/Q vssd1 vssd1 vccd1 vccd1 hold732/X sky130_fd_sc_hd__dlygate4sd3_1
X_1789_ _2121_/A _2059_/A vssd1 vssd1 vccd1 vccd1 _2123_/A sky130_fd_sc_hd__or2_1
X_3528_ _3542_/CLK _3528_/D _3022_/Y vssd1 vssd1 vccd1 vccd1 _3528_/Q sky130_fd_sc_hd__dfrtp_1
Xhold787 _2615_/X vssd1 vssd1 vccd1 vccd1 _3157_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 _3432_/Q vssd1 vssd1 vccd1 vccd1 hold776/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 _2851_/X vssd1 vssd1 vccd1 vccd1 _3374_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3459_ _3636_/CLK hold84/X _2953_/Y vssd1 vssd1 vccd1 vccd1 _3459_/Q sky130_fd_sc_hd__dfrtp_1
Xhold798 _3435_/Q vssd1 vssd1 vccd1 vccd1 hold798/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1961__S0 _1590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2761__S _2763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2594__A1 _2810_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2001__S _2045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold92 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_85_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2830_ hold580/X _2079_/A _2833_/S vssd1 vssd1 vccd1 vccd1 _2830_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2671__S _2672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2761_ hold390/X _2811_/A1 _2763_/S vssd1 vssd1 vccd1 vccd1 _2761_/X sky130_fd_sc_hd__mux2_1
X_1712_ _3531_/Q hold88/X vssd1 vssd1 vccd1 vccd1 _1712_/Y sky130_fd_sc_hd__nand2b_1
X_2692_ _2812_/A1 hold353/X _2693_/S vssd1 vssd1 vccd1 vccd1 _2692_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_1 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1643_ _2080_/A _2395_/A hold8/X vssd1 vssd1 vccd1 vccd1 _1643_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2432__S1 _1911_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1574_ _1574_/A vssd1 vssd1 vccd1 vccd1 _2350_/A sky130_fd_sc_hd__inv_2
X_3313_ _3488_/CLK _3313_/D vssd1 vssd1 vccd1 vccd1 _3313_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _3316_/CLK _3244_/D vssd1 vssd1 vccd1 vccd1 _3244_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3175_ _3583_/CLK _3175_/D vssd1 vssd1 vccd1 vccd1 _3175_/Q sky130_fd_sc_hd__dfxtp_1
X_2126_ _3502_/Q _2126_/B vssd1 vssd1 vccd1 vccd1 _2127_/D sky130_fd_sc_hd__xnor2_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2057_ _2054_/A _3625_/Q _2081_/C vssd1 vssd1 vccd1 vccd1 _2089_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_88_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2499__S1 _2550_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2959_ _3128_/A vssd1 vssd1 vccd1 vccd1 _2959_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2328__A1 _3443_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold551 _2818_/X vssd1 vssd1 vccd1 vccd1 _3335_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 _3356_/Q vssd1 vssd1 vccd1 vccd1 hold562/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold540 _3338_/Q vssd1 vssd1 vccd1 vccd1 hold540/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 _2654_/X vssd1 vssd1 vccd1 vccd1 _3190_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 _3189_/Q vssd1 vssd1 vccd1 vccd1 hold584/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 _2873_/X vssd1 vssd1 vccd1 vccd1 _3399_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2756__S _2763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput60 _3659_/A vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_12
XANTENNA__2666__S _2672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2813_ hold418/X _2813_/A1 _2813_/S vssd1 vssd1 vccd1 vccd1 _2813_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2744_ _2784_/C _2794_/A _2794_/B vssd1 vssd1 vccd1 vccd1 _2753_/S sky130_fd_sc_hd__or3b_4
X_2675_ hold169/X _2806_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2675_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1626_ _1626_/A vssd1 vssd1 vccd1 vccd1 _1668_/A sky130_fd_sc_hd__inv_2
X_1557_ _1557_/A vssd1 vssd1 vccd1 vccd1 _1692_/A sky130_fd_sc_hd__inv_2
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3227_ _3328_/CLK _3227_/D vssd1 vssd1 vccd1 vccd1 _3227_/Q sky130_fd_sc_hd__dfxtp_1
X_3158_ _3416_/CLK _3158_/D vssd1 vssd1 vccd1 vccd1 _3158_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2494__A0 _3341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2109_ _2108_/A _2081_/B _2108_/Y _2076_/B vssd1 vssd1 vccd1 vccd1 _2109_/X sky130_fd_sc_hd__o211a_2
X_3089_ _3089_/A vssd1 vssd1 vccd1 vccd1 _3089_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_49_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2797__A1 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold381 _2753_/X vssd1 vssd1 vccd1 vccd1 _3277_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold370 _3221_/Q vssd1 vssd1 vccd1 vccd1 hold370/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 _3255_/Q vssd1 vssd1 vccd1 vccd1 hold392/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2486__S _2551_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3319_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2460_ _3485_/Q _2507_/C _2508_/A vssd1 vssd1 vccd1 vccd1 _2460_/X sky130_fd_sc_hd__o21a_1
X_2391_ _2391_/A _2391_/B _2391_/C vssd1 vssd1 vccd1 vccd1 _2391_/X sky130_fd_sc_hd__or3_2
XFILLER_0_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3012_ _3114_/A vssd1 vssd1 vccd1 vccd1 _3012_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_6_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout127_A _3131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2727_ _2807_/A1 hold272/X _2733_/S vssd1 vssd1 vccd1 vccd1 _2727_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2658_ _2075_/B hold732/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2658_/X sky130_fd_sc_hd__mux2_1
Xfanout113 hold176/X vssd1 vssd1 vccd1 vccd1 _2585_/A sky130_fd_sc_hd__clkbuf_4
X_1609_ _1609_/A _1609_/B _1907_/B vssd1 vssd1 vccd1 vccd1 _2393_/A sky130_fd_sc_hd__nand3_4
Xfanout102 hold44/X vssd1 vssd1 vccd1 vccd1 _2812_/A1 sky130_fd_sc_hd__clkbuf_4
X_2589_ hold360/X _2805_/A1 _2594_/S vssd1 vssd1 vccd1 vccd1 _2589_/X sky130_fd_sc_hd__mux2_1
Xfanout124 _3089_/A vssd1 vssd1 vccd1 vccd1 _3126_/A sky130_fd_sc_hd__buf_8
XFILLER_0_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1690__A1 _2585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2553__S0 _2554_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1681__A1 hold14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1960_ _1958_/X _1959_/X _2045_/S vssd1 vssd1 vccd1 vccd1 _1960_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1891_ _1891_/A _2231_/D vssd1 vssd1 vccd1 vccd1 _2630_/C sky130_fd_sc_hd__or2_2
XFILLER_0_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3630_ _3631_/CLK hold91/X _3121_/Y vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__dfrtp_1
X_3561_ _3563_/CLK _3561_/D _3055_/Y vssd1 vssd1 vccd1 vccd1 _3561_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_51_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2512_ hold79/A _2568_/B _2417_/B _3377_/Q _2509_/X vssd1 vssd1 vccd1 vccd1 _2512_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3492_ _3493_/CLK _3492_/D _2986_/Y vssd1 vssd1 vccd1 vccd1 _3492_/Q sky130_fd_sc_hd__dfrtp_4
X_2443_ _2440_/X _2508_/B _2442_/X _2441_/A _3608_/Q vssd1 vssd1 vccd1 vccd1 _2443_/X
+ sky130_fd_sc_hd__a32o_1
X_2374_ _1824_/A _1793_/A _2370_/Y _2373_/X vssd1 vssd1 vccd1 vccd1 _2374_/X sky130_fd_sc_hd__a31o_1
XANTENNA__2697__A0 _2807_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2544__S0 _2554_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2621__A0 _2342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2688__A0 _2808_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2860__A0 _2111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2612__A0 _2105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2004__S _2045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output40_A _3581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2090_ _2121_/A _3546_/Q _2089_/B _2088_/Y vssd1 vssd1 vccd1 vccd1 _2090_/X sky130_fd_sc_hd__a31o_1
XANTENNA__2674__S _2682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1654__A1 _2396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2992_ _3065_/A vssd1 vssd1 vccd1 vccd1 _2992_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_83_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2603__A0 _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1943_ _3523_/Q _1943_/B vssd1 vssd1 vccd1 vccd1 _1944_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1874_ _1873_/Y _1871_/B _1843_/A _1560_/Y vssd1 vssd1 vccd1 vccd1 _3533_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3613_ _3614_/CLK _3613_/D _3104_/Y vssd1 vssd1 vccd1 vccd1 _3613_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_hold65_A hold65/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold903 _1705_/Y vssd1 vssd1 vccd1 vccd1 hold903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 _1876_/X vssd1 vssd1 vccd1 vccd1 _3532_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3544_ _3583_/CLK _3544_/D _3038_/Y vssd1 vssd1 vccd1 vccd1 _3544_/Q sky130_fd_sc_hd__dfrtp_1
Xhold914 _1707_/B vssd1 vssd1 vccd1 vccd1 hold914/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 _3571_/Q vssd1 vssd1 vccd1 vccd1 hold925/X sky130_fd_sc_hd__dlygate4sd3_1
X_3475_ _3583_/CLK _3475_/D _2969_/Y vssd1 vssd1 vccd1 vccd1 _3475_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold947 _1902_/Y vssd1 vssd1 vccd1 vccd1 hold947/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 _1773_/X vssd1 vssd1 vccd1 vccd1 _3560_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 _3563_/Q vssd1 vssd1 vccd1 vccd1 _1761_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2426_ _3638_/Q _2511_/A _2405_/Y _2425_/X vssd1 vssd1 vccd1 vccd1 _2426_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_86_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2357_ _1577_/Y _2208_/A _2205_/A _1578_/Y _2356_/X vssd1 vssd1 vccd1 vccd1 _2357_/X
+ sky130_fd_sc_hd__a221o_1
X_2288_ hold18/X _2409_/B vssd1 vssd1 vccd1 vccd1 _2419_/B sky130_fd_sc_hd__nor2_2
XANTENNA__2842__A0 _2338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2759__S _2763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1636__A1 hold49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1590_ _1590_/A vssd1 vssd1 vccd1 vccd1 _2196_/A sky130_fd_sc_hd__inv_2
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2669__S _2672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _3305_/CLK _3260_/D vssd1 vssd1 vccd1 vccd1 _3260_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ _2211_/A _2211_/B vssd1 vssd1 vccd1 vccd1 _2211_/X sky130_fd_sc_hd__xor2_1
X_3191_ _3403_/CLK _3191_/D vssd1 vssd1 vccd1 vccd1 _3191_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2142_ _2136_/C _2141_/X hold962/X vssd1 vssd1 vccd1 vccd1 _2142_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2073_ _2080_/A _2070_/X _2072_/Y vssd1 vssd1 vccd1 vccd1 _2073_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_88_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2052__A1 _2320_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2975_ _3065_/A vssd1 vssd1 vccd1 vccd1 _2975_/Y sky130_fd_sc_hd__inv_2
X_1926_ _1940_/S _1938_/B vssd1 vssd1 vccd1 vccd1 _1926_/Y sky130_fd_sc_hd__nand2_1
X_1857_ _1859_/A _1835_/A _1859_/B _1853_/A vssd1 vssd1 vccd1 vccd1 _1858_/B sky130_fd_sc_hd__a31o_1
Xhold700 _3361_/Q vssd1 vssd1 vccd1 vccd1 hold700/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold711 _2600_/X vssd1 vssd1 vccd1 vccd1 _3143_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3527_ _3542_/CLK _3527_/D _3021_/Y vssd1 vssd1 vccd1 vccd1 _3527_/Q sky130_fd_sc_hd__dfrtp_2
Xhold755 _2605_/X vssd1 vssd1 vccd1 vccd1 _3148_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 _3430_/Q vssd1 vssd1 vccd1 vccd1 hold744/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 _3404_/Q vssd1 vssd1 vccd1 vccd1 hold722/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 _2658_/X vssd1 vssd1 vccd1 vccd1 _3194_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1788_ _3627_/Q _2056_/A vssd1 vssd1 vccd1 vccd1 _2059_/A sky130_fd_sc_hd__or2_2
XFILLER_0_12_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold766 _3150_/Q vssd1 vssd1 vccd1 vccd1 hold766/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 _2910_/X vssd1 vssd1 vccd1 vccd1 _3432_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold788 _3144_/Q vssd1 vssd1 vccd1 vccd1 hold788/X sky130_fd_sc_hd__dlygate4sd3_1
X_3458_ _3636_/CLK hold12/X _2952_/Y vssd1 vssd1 vccd1 vccd1 _3458_/Q sky130_fd_sc_hd__dfrtp_1
Xhold799 _2913_/X vssd1 vssd1 vccd1 vccd1 _3435_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3389_ _3436_/CLK _3389_/D vssd1 vssd1 vccd1 vccd1 _3389_/Q sky130_fd_sc_hd__dfxtp_1
X_2409_ _2418_/B _2409_/B vssd1 vssd1 vccd1 vccd1 _2441_/B sky130_fd_sc_hd__nor2_1
XANTENNA__1961__S1 _2193_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3579_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold82 wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__buf_2
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2760_ hold343/X _2810_/A1 _2763_/S vssd1 vssd1 vccd1 vccd1 _2760_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1711_ _1711_/A _1711_/B vssd1 vssd1 vccd1 vccd1 _1711_/X sky130_fd_sc_hd__xor2_1
X_2691_ _2811_/A1 hold370/X _2693_/S vssd1 vssd1 vccd1 vccd1 _2691_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1642_ _2054_/A _2396_/A hold8/X vssd1 vssd1 vccd1 vccd1 _1642_/X sky130_fd_sc_hd__mux2_1
XANTENNA_2 hold44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1573_ _1573_/A vssd1 vssd1 vccd1 vccd1 _1573_/Y sky130_fd_sc_hd__inv_2
X_3312_ _3488_/CLK _3312_/D vssd1 vssd1 vccd1 vccd1 _3312_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _3319_/CLK _3243_/D vssd1 vssd1 vccd1 vccd1 _3243_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ _3423_/CLK _3174_/D vssd1 vssd1 vccd1 vccd1 _3174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2125_ _2125_/A _2321_/B vssd1 vssd1 vccd1 vccd1 _2127_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2056_ _2056_/A _2056_/B vssd1 vssd1 vccd1 vccd1 _2108_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_76_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2862__S _2864_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2958_ _3128_/A vssd1 vssd1 vccd1 vccd1 _2958_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1909_ _1933_/A _1909_/B vssd1 vssd1 vccd1 vccd1 _1910_/B sky130_fd_sc_hd__nor2_2
X_2889_ _2104_/X hold646/X _2894_/S vssd1 vssd1 vccd1 vccd1 _2889_/X sky130_fd_sc_hd__mux2_1
Xhold530 _3427_/Q vssd1 vssd1 vccd1 vccd1 hold530/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 _3333_/Q vssd1 vssd1 vccd1 vccd1 hold552/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 _2831_/X vssd1 vssd1 vccd1 vccd1 _3356_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold541 _2821_/X vssd1 vssd1 vccd1 vccd1 _3338_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 _3193_/Q vssd1 vssd1 vccd1 vccd1 hold596/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 _2653_/X vssd1 vssd1 vccd1 vccd1 _3189_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 _3178_/Q vssd1 vssd1 vccd1 vccd1 hold574/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2772__S _2773_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput61 _2491_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_12
Xoutput50 _3652_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_12
XANTENNA__2012__S _2045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2682__S _2682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2812_ hold382/X _2812_/A1 _2813_/S vssd1 vssd1 vccd1 vccd1 _2812_/X sky130_fd_sc_hd__mux2_1
X_2743_ _2813_/A1 hold347/X _2743_/S vssd1 vssd1 vccd1 vccd1 _2743_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2674_ hold261/X _2805_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2674_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1625_ hold93/X _1625_/B hold17/X _1613_/B vssd1 vssd1 vccd1 vccd1 _1625_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_1_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2857__S _2864_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3226_ _3325_/CLK _3226_/D vssd1 vssd1 vccd1 vccd1 _3226_/Q sky130_fd_sc_hd__dfxtp_1
X_3157_ _3583_/CLK _3157_/D vssd1 vssd1 vccd1 vccd1 _3157_/Q sky130_fd_sc_hd__dfxtp_1
X_2108_ _2108_/A _2108_/B vssd1 vssd1 vccd1 vccd1 _2108_/Y sky130_fd_sc_hd__nand2_1
X_3088_ _3124_/A vssd1 vssd1 vccd1 vccd1 _3088_/Y sky130_fd_sc_hd__inv_2
X_2039_ _1985_/S _2034_/X _2038_/X vssd1 vssd1 vccd1 vccd1 _2039_/Y sky130_fd_sc_hd__a21oi_2
Xhold371 _2691_/X vssd1 vssd1 vccd1 vccd1 _3221_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold360 _3134_/Q vssd1 vssd1 vccd1 vccd1 hold360/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2767__S _2773_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold393 _2729_/X vssd1 vssd1 vccd1 vccd1 _3255_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _3330_/Q vssd1 vssd1 vccd1 vccd1 hold382/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1060 _3517_/Q vssd1 vssd1 vccd1 vccd1 hold500/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2390_ _3597_/Q _3382_/Q _3341_/Q _3600_/Q _2388_/X vssd1 vssd1 vccd1 vccd1 _2391_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2677__S _2682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3011_ _3114_/A vssd1 vssd1 vccd1 vccd1 _3011_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1610__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2726_ _2806_/A1 hold191/X _2733_/S vssd1 vssd1 vccd1 vccd1 _2726_/X sky130_fd_sc_hd__mux2_1
X_2657_ _2079_/A hold596/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2657_/X sky130_fd_sc_hd__mux2_1
X_1608_ _1609_/A _1609_/B _1907_/B vssd1 vssd1 vccd1 vccd1 _2585_/B sky130_fd_sc_hd__and3_1
Xfanout103 hold52/X vssd1 vssd1 vccd1 vccd1 _2811_/A1 sky130_fd_sc_hd__clkbuf_4
X_2588_ _2794_/B _2794_/C _2794_/A vssd1 vssd1 vccd1 vccd1 _2597_/S sky130_fd_sc_hd__nor3b_4
Xfanout125 _3131_/A vssd1 vssd1 vccd1 vccd1 _3133_/A sky130_fd_sc_hd__buf_8
XFILLER_0_10_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout114 _3120_/A vssd1 vssd1 vccd1 vccd1 _3114_/A sky130_fd_sc_hd__buf_8
XANTENNA__2011__S0 _2044_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3209_ _3328_/CLK _3209_/D vssd1 vssd1 vccd1 vccd1 _3209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold190 _2756_/X vssd1 vssd1 vccd1 vccd1 _3279_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2002__S0 _2044_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2553__S1 _1911_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1890_ _1891_/A _2231_/D vssd1 vssd1 vccd1 vccd1 _2598_/C sky130_fd_sc_hd__nor2_4
XFILLER_0_50_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3560_ _3563_/CLK _3560_/D _3054_/Y vssd1 vssd1 vccd1 vccd1 _3560_/Q sky130_fd_sc_hd__dfstp_1
X_2511_ _2511_/A _2511_/B vssd1 vssd1 vccd1 vccd1 _2511_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_59_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3491_ _3493_/CLK _3491_/D _2985_/Y vssd1 vssd1 vccd1 vccd1 _3491_/Q sky130_fd_sc_hd__dfrtp_4
X_2442_ _3597_/Q _2568_/B vssd1 vssd1 vccd1 vccd1 _2442_/X sky130_fd_sc_hd__or2_1
X_2373_ _1808_/B _1808_/D _2383_/C vssd1 vssd1 vccd1 vccd1 _2373_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2544__S1 _1911_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2709_ _2809_/A1 hold410/X _2713_/S vssd1 vssd1 vccd1 vccd1 _2709_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2231__D _2231_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2679__A1 _2810_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2020__S _2053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2690__S _2693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2991_ _3131_/A vssd1 vssd1 vccd1 vccd1 _2991_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1942_ _1942_/A _1942_/B vssd1 vssd1 vccd1 vccd1 _2165_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1873_ _1843_/A _1843_/B _1835_/A vssd1 vssd1 vccd1 vccd1 _1873_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3087__A _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3612_ _3612_/CLK _3612_/D _3103_/Y vssd1 vssd1 vccd1 vccd1 _3612_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold904 _1706_/Y vssd1 vssd1 vccd1 vccd1 _3575_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold915 _3540_/Q vssd1 vssd1 vccd1 vccd1 _1859_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3543_ _3583_/CLK _3543_/D _3037_/Y vssd1 vssd1 vccd1 vccd1 _3543_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold937 _3642_/Q vssd1 vssd1 vccd1 vccd1 _1557_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 _1748_/X vssd1 vssd1 vccd1 vccd1 _3571_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3474_ _3583_/CLK _3474_/D _2968_/Y vssd1 vssd1 vccd1 vccd1 _3474_/Q sky130_fd_sc_hd__dfrtp_1
Xhold959 _3525_/Q vssd1 vssd1 vccd1 vccd1 hold959/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold948 _1903_/Y vssd1 vssd1 vccd1 vccd1 _3524_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_2_2__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2425_ _3615_/Q _1645_/Y _2408_/X _2424_/X vssd1 vssd1 vccd1 vccd1 _2425_/X sky130_fd_sc_hd__a22o_1
X_2356_ _1578_/Y _2205_/A _2220_/S _1579_/Y vssd1 vssd1 vccd1 vccd1 _2356_/X sky130_fd_sc_hd__o22a_1
X_2287_ _2287_/A hold57/X hold5/X _1657_/C vssd1 vssd1 vccd1 vccd1 _2287_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_79_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2833__A1 _2339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2015__S _2045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _2207_/A _2207_/B _2216_/B vssd1 vssd1 vccd1 vccd1 _2212_/B sky130_fd_sc_hd__a21bo_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _3369_/CLK _3190_/D vssd1 vssd1 vccd1 vccd1 _3190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2141_ _2134_/B _2134_/C _2052_/S vssd1 vssd1 vccd1 vccd1 _2141_/X sky130_fd_sc_hd__a21o_1
XANTENNA__2685__S _2693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2072_ _2080_/A _2080_/B vssd1 vssd1 vccd1 vccd1 _2072_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2974_ _3065_/A vssd1 vssd1 vccd1 vccd1 _2974_/Y sky130_fd_sc_hd__inv_2
X_1925_ _2350_/B _1931_/B vssd1 vssd1 vccd1 vccd1 _1938_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_44_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_6_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3612_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1856_ _1855_/A _1858_/A _1855_/Y _1853_/X vssd1 vssd1 vccd1 vccd1 _1856_/X sky130_fd_sc_hd__a22o_1
Xhold701 _2837_/X vssd1 vssd1 vccd1 vccd1 _3361_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 _3145_/Q vssd1 vssd1 vccd1 vccd1 hold712/X sky130_fd_sc_hd__dlygate4sd3_1
X_1787_ _2121_/A _3556_/Q vssd1 vssd1 vccd1 vccd1 _1787_/X sky130_fd_sc_hd__or2_1
XFILLER_0_52_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold723 _2879_/X vssd1 vssd1 vccd1 vccd1 _3404_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold734 _3186_/Q vssd1 vssd1 vccd1 vccd1 hold734/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 _2908_/X vssd1 vssd1 vccd1 vccd1 _3430_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3526_ _3526_/CLK _3526_/D _3020_/Y vssd1 vssd1 vccd1 vccd1 _3526_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout102_A hold44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold778 _3375_/Q vssd1 vssd1 vccd1 vccd1 hold778/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 _2607_/X vssd1 vssd1 vccd1 vccd1 _3150_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 _3384_/Q vssd1 vssd1 vccd1 vccd1 hold756/X sky130_fd_sc_hd__dlygate4sd3_1
X_3457_ _3637_/CLK hold37/X _2951_/Y vssd1 vssd1 vccd1 vccd1 _3457_/Q sky130_fd_sc_hd__dfrtp_1
Xhold789 _2601_/X vssd1 vssd1 vccd1 vccd1 _3144_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3388_ _3433_/CLK _3388_/D vssd1 vssd1 vccd1 vccd1 _3388_/Q sky130_fd_sc_hd__dfxtp_1
X_2408_ _3515_/Q _2507_/B hold59/A vssd1 vssd1 vccd1 vccd1 _2408_/X sky130_fd_sc_hd__o21a_1
X_2339_ _3623_/Q _2339_/B vssd1 vssd1 vccd1 vccd1 _2339_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2815__A1 _2342_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2751__A0 _2811_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__buf_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2806__A1 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1710_ hold914/X _1709_/Y _3466_/D vssd1 vssd1 vccd1 vccd1 _3573_/D sky130_fd_sc_hd__a21oi_1
X_2690_ _2810_/A1 hold302/X _2693_/S vssd1 vssd1 vccd1 vccd1 _2690_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_3 _2339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1641_ _2081_/C _2397_/A hold8/X vssd1 vssd1 vccd1 vccd1 _1641_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2742__A0 _2812_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3311_ _3488_/CLK _3311_/D vssd1 vssd1 vccd1 vccd1 _3311_/Q sky130_fd_sc_hd__dfxtp_1
X_1572_ _3614_/Q vssd1 vssd1 vccd1 vccd1 _1572_/Y sky130_fd_sc_hd__inv_2
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ _3316_/CLK _3242_/D vssd1 vssd1 vccd1 vccd1 _3242_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ _3369_/CLK _3173_/D vssd1 vssd1 vccd1 vccd1 _3173_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2124_ _2134_/B _2124_/B vssd1 vssd1 vccd1 vccd1 _2127_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_83_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2055_ _2056_/A _2056_/B vssd1 vssd1 vccd1 vccd1 _2082_/A sky130_fd_sc_hd__and2_1
X_2957_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2957_/Y sky130_fd_sc_hd__inv_2
X_2888_ _2101_/X hold636/X _2894_/S vssd1 vssd1 vccd1 vccd1 _2888_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1908_ _1921_/A _2630_/C _1922_/B vssd1 vssd1 vccd1 vccd1 _1909_/B sky130_fd_sc_hd__a21oi_1
X_1839_ _1877_/B vssd1 vssd1 vccd1 vccd1 _1839_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold520 _3358_/Q vssd1 vssd1 vccd1 vccd1 hold520/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 _2816_/X vssd1 vssd1 vccd1 vccd1 _3333_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 _3334_/Q vssd1 vssd1 vccd1 vccd1 hold542/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 _2904_/X vssd1 vssd1 vccd1 vccd1 _3427_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2733__A0 _2813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold586 _3415_/Q vssd1 vssd1 vccd1 vccd1 hold586/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 _2657_/X vssd1 vssd1 vccd1 vccd1 _3193_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 _3423_/Q vssd1 vssd1 vccd1 vccd1 hold564/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold575 _2640_/X vssd1 vssd1 vccd1 vccd1 _3178_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3509_ _3513_/CLK _3509_/D _3003_/Y vssd1 vssd1 vccd1 vccd1 _3509_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2338__B _2338_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput40 _3581_/Q vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_12
Xoutput51 _2455_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_12
XFILLER_0_31_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput62 _2506_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_12
XFILLER_0_73_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2811_ hold412/X _2811_/A1 _2813_/S vssd1 vssd1 vccd1 vccd1 _2811_/X sky130_fd_sc_hd__mux2_1
X_2742_ _2812_/A1 hold313/X _2743_/S vssd1 vssd1 vccd1 vccd1 _2742_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_82_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1608__A _1609_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2673_ _2794_/C _2804_/B vssd1 vssd1 vccd1 vccd1 _2682_/S sky130_fd_sc_hd__nor2_4
XANTENNA__2715__A0 _2805_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1624_ _2287_/A input3/X _1624_/C hold5/X vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__or4_2
X_3225_ _3328_/CLK _3225_/D vssd1 vssd1 vccd1 vccd1 _3225_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3156_ _3414_/CLK _3156_/D vssd1 vssd1 vccd1 vccd1 _3156_/Q sky130_fd_sc_hd__dfxtp_1
X_3087_ _3089_/A vssd1 vssd1 vccd1 vccd1 _3087_/Y sky130_fd_sc_hd__inv_2
X_2107_ _2107_/A _2107_/B vssd1 vssd1 vccd1 vccd1 _2112_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2038_ _1985_/S _2038_/B vssd1 vssd1 vccd1 vccd1 _2038_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_64_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2706__A0 _2806_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold350 _2793_/X vssd1 vssd1 vccd1 vccd1 _3313_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 _2589_/X vssd1 vssd1 vccd1 vccd1 _3134_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 _3311_/Q vssd1 vssd1 vccd1 vccd1 hold372/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 _3230_/Q vssd1 vssd1 vccd1 vccd1 hold394/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 _2812_/X vssd1 vssd1 vccd1 vccd1 _3330_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1050 wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2023__S _2045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3633_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1920__A1 _1911_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3010_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3010_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2693__S _2693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1610__B input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2725_ _2805_/A1 hold307/X _2733_/S vssd1 vssd1 vccd1 vccd1 _2725_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2656_ _2111_/B hold662/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2656_/X sky130_fd_sc_hd__mux2_1
X_1607_ _1609_/A _1609_/B vssd1 vssd1 vccd1 vccd1 _2586_/B sky130_fd_sc_hd__nand2_1
Xfanout104 hold33/X vssd1 vssd1 vccd1 vccd1 _2810_/A1 sky130_fd_sc_hd__buf_4
X_2587_ _3492_/Q _3491_/Q _2587_/C vssd1 vssd1 vccd1 vccd1 _2794_/C sky130_fd_sc_hd__nand3b_4
Xfanout115 _3089_/A vssd1 vssd1 vccd1 vccd1 _3120_/A sky130_fd_sc_hd__buf_6
Xfanout126 _3131_/A vssd1 vssd1 vccd1 vccd1 _3065_/A sky130_fd_sc_hd__buf_8
X_3208_ _3325_/CLK _3208_/D vssd1 vssd1 vccd1 vccd1 _3208_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1675__A0 _2585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2011__S1 _2044_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3139_ _3330_/CLK _3139_/D vssd1 vssd1 vccd1 vccd1 _3139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold180 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 input19/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 _3252_/Q vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2079__A _2079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2002__S1 _2044_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3490_ _3610_/CLK _3490_/D _2984_/Y vssd1 vssd1 vccd1 vccd1 _3490_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2510_ hold80/A hold7/A vssd1 vssd1 vccd1 vccd1 _2510_/X sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2688__S _2693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2441_ _2441_/A _2441_/B vssd1 vssd1 vccd1 vccd1 _2508_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2372_ _2371_/X _2378_/B _2379_/S vssd1 vssd1 vccd1 vccd1 _2372_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2909__A0 _2105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2708_ _2808_/A1 hold134/X _2713_/S vssd1 vssd1 vccd1 vccd1 _2708_/X sky130_fd_sc_hd__mux2_1
X_2639_ _2338_/B hold758/X _2640_/S vssd1 vssd1 vccd1 vccd1 _2639_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1991__S0 _1590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1982__S0 _1590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2300__A1 hold44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2990_ _3065_/A vssd1 vssd1 vccd1 vccd1 _2990_/Y sky130_fd_sc_hd__inv_2
X_1941_ _3524_/Q _3523_/Q vssd1 vssd1 vccd1 vccd1 _1942_/B sky130_fd_sc_hd__xor2_1
X_1872_ _1835_/A _1844_/Y _1871_/X _1871_/A _1560_/Y vssd1 vssd1 vccd1 vccd1 _1872_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3611_ _3612_/CLK _3611_/D _3102_/Y vssd1 vssd1 vccd1 vccd1 _3611_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold916 _1860_/X vssd1 vssd1 vccd1 vccd1 _3540_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3542_ _3542_/CLK _3542_/D _3036_/Y vssd1 vssd1 vccd1 vccd1 _3542_/Q sky130_fd_sc_hd__dfrtp_1
Xhold905 _3442_/Q vssd1 vssd1 vccd1 vccd1 _1808_/D sky130_fd_sc_hd__buf_1
Xhold927 _3437_/Q vssd1 vssd1 vccd1 vccd1 hold927/X sky130_fd_sc_hd__dlygate4sd3_1
X_3473_ _3576_/CLK _3473_/D _2967_/Y vssd1 vssd1 vccd1 vccd1 _3473_/Q sky130_fd_sc_hd__dfrtp_1
Xhold949 _3569_/Q vssd1 vssd1 vccd1 vccd1 _1749_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold938 _3497_/Q vssd1 vssd1 vccd1 vccd1 _2129_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2424_ _2423_/X _3611_/Q _2439_/A vssd1 vssd1 vccd1 vccd1 _2424_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2355_ _2353_/X _2354_/X hold909/X vssd1 vssd1 vccd1 vccd1 _2355_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_19_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2286_ _2272_/B _2272_/C _2285_/Y vssd1 vssd1 vccd1 vccd1 _2286_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_79_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1960__S _2045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2791__S _2793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2092__A _2097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2597__A1 _2813_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2031__S _2053_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3651__A _3659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2140_ _2134_/C _2136_/C _2134_/B vssd1 vssd1 vccd1 vccd1 _2140_/Y sky130_fd_sc_hd__a21oi_1
X_2071_ _2071_/A _2071_/B vssd1 vssd1 vccd1 vccd1 _2080_/B sky130_fd_sc_hd__or2_2
XFILLER_0_88_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2973_ _3065_/A vssd1 vssd1 vccd1 vccd1 _2973_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3098__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1924_ _1928_/A _1931_/B vssd1 vssd1 vccd1 vccd1 _1929_/A sky130_fd_sc_hd__and2_1
XFILLER_0_16_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1855_ _1855_/A _1855_/B vssd1 vssd1 vccd1 vccd1 _1855_/Y sky130_fd_sc_hd__nor2_1
Xhold702 _3360_/Q vssd1 vssd1 vccd1 vccd1 hold702/X sky130_fd_sc_hd__dlygate4sd3_1
X_1786_ _2121_/A _3556_/Q vssd1 vssd1 vccd1 vccd1 _1786_/Y sky130_fd_sc_hd__nand2_1
Xhold746 _3366_/Q vssd1 vssd1 vccd1 vccd1 hold746/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 _2649_/X vssd1 vssd1 vccd1 vccd1 _3186_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 _2602_/X vssd1 vssd1 vccd1 vccd1 _3145_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 _3363_/Q vssd1 vssd1 vccd1 vccd1 hold724/X sky130_fd_sc_hd__dlygate4sd3_1
X_3525_ _3526_/CLK _3525_/D _3019_/Y vssd1 vssd1 vccd1 vccd1 _3525_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__2760__A1 _2810_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold779 _2852_/X vssd1 vssd1 vccd1 vccd1 _3375_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 _2857_/X vssd1 vssd1 vccd1 vccd1 _3384_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 _3405_/Q vssd1 vssd1 vccd1 vccd1 hold768/X sky130_fd_sc_hd__dlygate4sd3_1
X_3456_ _3540_/CLK hold77/X _2950_/Y vssd1 vssd1 vccd1 vccd1 _3456_/Q sky130_fd_sc_hd__dfrtp_1
X_3387_ _3404_/CLK _3387_/D vssd1 vssd1 vccd1 vccd1 _3387_/Q sky130_fd_sc_hd__dfxtp_1
X_2407_ _2407_/A hold19/A vssd1 vssd1 vccd1 vccd1 _2507_/B sky130_fd_sc_hd__nand2_1
X_2338_ hold69/A _2338_/B vssd1 vssd1 vccd1 vccd1 _2338_/Y sky130_fd_sc_hd__xnor2_1
X_2269_ _2268_/X _2269_/B _2269_/C _2269_/D vssd1 vssd1 vccd1 vccd1 _2269_/X sky130_fd_sc_hd__and4b_1
XFILLER_0_67_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2786__S _2793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_45_wb_clk_i clkbuf_leaf_5_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3423_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2026__S _2045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1640_ _2383_/A hold86/X hold8/X vssd1 vssd1 vccd1 vccd1 _1640_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1571_ _1571_/A vssd1 vssd1 vccd1 vccd1 _1571_/Y sky130_fd_sc_hd__inv_2
X_3310_ _3319_/CLK _3310_/D vssd1 vssd1 vccd1 vccd1 _3310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _3513_/CLK _3241_/D vssd1 vssd1 vccd1 vccd1 _3241_/Q sky130_fd_sc_hd__dfxtp_1
X_3172_ _3582_/CLK _3172_/D vssd1 vssd1 vccd1 vccd1 _3172_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2123_ _2123_/A _2123_/B _2123_/C vssd1 vssd1 vccd1 vccd1 _2127_/A sky130_fd_sc_hd__and3_1
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2054_ _2054_/A _3625_/Q vssd1 vssd1 vccd1 vccd1 _2056_/B sky130_fd_sc_hd__nand2_2
X_2956_ _3124_/A vssd1 vssd1 vccd1 vccd1 _2956_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2887_ _2091_/X hold652/X _2894_/S vssd1 vssd1 vccd1 vccd1 _2887_/X sky130_fd_sc_hd__mux2_1
X_1907_ _2586_/B _1907_/B _3581_/Q _2506_/S vssd1 vssd1 vccd1 vccd1 _1922_/B sky130_fd_sc_hd__or4bb_4
XFILLER_0_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1838_ _1838_/A _1838_/B _3528_/Q _3527_/Q vssd1 vssd1 vccd1 vccd1 _1877_/B sky130_fd_sc_hd__and4_2
XFILLER_0_4_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold510 _3592_/Q vssd1 vssd1 vccd1 vccd1 _2333_/A sky130_fd_sc_hd__dlygate4sd3_1
X_1769_ hold826/X _3475_/Q _3642_/Q vssd1 vssd1 vccd1 vccd1 _1769_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold532 _3352_/Q vssd1 vssd1 vccd1 vccd1 hold532/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 _2817_/X vssd1 vssd1 vccd1 vccd1 _3334_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 _3332_/Q vssd1 vssd1 vccd1 vccd1 hold554/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold521 _2833_/X vssd1 vssd1 vccd1 vccd1 _3358_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 _2891_/X vssd1 vssd1 vccd1 vccd1 _3415_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold576 _3421_/Q vssd1 vssd1 vccd1 vccd1 hold576/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 _2900_/X vssd1 vssd1 vccd1 vccd1 _3423_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3508_ _3513_/CLK _3508_/D _3002_/Y vssd1 vssd1 vccd1 vccd1 _3508_/Q sky130_fd_sc_hd__dfrtp_1
Xhold598 _3433_/Q vssd1 vssd1 vccd1 vccd1 hold598/X sky130_fd_sc_hd__dlygate4sd3_1
X_3439_ _3559_/CLK _3439_/D _2933_/Y vssd1 vssd1 vccd1 vccd1 _3439_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput52 _3653_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_12
Xoutput41 _2435_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_12
Xoutput63 _2522_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_12
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2660__A0 _2339_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2810_ hold351/X _2810_/A1 _2813_/S vssd1 vssd1 vccd1 vccd1 _2810_/X sky130_fd_sc_hd__mux2_1
X_2741_ _2811_/A1 hold333/X _2743_/S vssd1 vssd1 vccd1 vccd1 _2741_/X sky130_fd_sc_hd__mux2_1
X_2672_ _2813_/A1 hold404/X _2672_/S vssd1 vssd1 vccd1 vccd1 _2672_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1608__B _1609_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1623_ _1834_/A _2585_/A _1623_/S vssd1 vssd1 vccd1 vccd1 _3638_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1624__A _2287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3224_ _3330_/CLK _3224_/D vssd1 vssd1 vccd1 vccd1 _3224_/Q sky130_fd_sc_hd__dfxtp_1
.ends

